
module Cipher ( clk, rst, Input, Key, Output );
  input [15:0] Input;
  input [31:0] Key;
  output [15:0] Output;
  (* SILVER="clock" *)input clk; 
  (* SILVER="control" *)input rst; 
  wire   AddKeyXOR1_XORInst_0_0_n1, AddKeyXOR1_XORInst_0_1_n1,
         AddKeyXOR1_XORInst_0_2_n1, AddKeyXOR1_XORInst_0_3_n1,
         AddKeyXOR1_XORInst_1_0_n1, AddKeyXOR1_XORInst_1_1_n1,
         AddKeyXOR1_XORInst_1_2_n1, AddKeyXOR1_XORInst_1_3_n1,
         AddKeyXOR1_XORInst_2_0_n1, AddKeyXOR1_XORInst_2_1_n1,
         AddKeyXOR1_XORInst_2_2_n1, AddKeyXOR1_XORInst_2_3_n1,
         AddKeyXOR1_XORInst_3_0_n1, AddKeyXOR1_XORInst_3_1_n1,
         AddKeyXOR1_XORInst_3_2_n1, AddKeyXOR1_XORInst_3_3_n1,
         AddKeyXOR2_XORInst_0_0_n1, AddKeyXOR2_XORInst_0_1_n1,
         AddKeyXOR2_XORInst_0_2_n1, AddKeyXOR2_XORInst_0_3_n1,
         AddKeyXOR2_XORInst_1_0_n1, AddKeyXOR2_XORInst_1_1_n1,
         AddKeyXOR2_XORInst_1_2_n1, AddKeyXOR2_XORInst_1_3_n1,
         AddKeyXOR2_XORInst_2_0_n1, AddKeyXOR2_XORInst_2_1_n1,
         AddKeyXOR2_XORInst_2_2_n1, AddKeyXOR2_XORInst_2_3_n1,
         AddKeyXOR2_XORInst_3_0_n1, AddKeyXOR2_XORInst_3_1_n1,
         AddKeyXOR2_XORInst_3_2_n1, AddKeyXOR2_XORInst_3_3_n1, n165, n166,
         n167, n168, n171, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360;

  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(AddKeyXOR1_XORInst_0_0_n1), .CK(
        clk), .Q(n197), .QN(n196) );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(AddKeyXOR1_XORInst_0_1_n1), .CK(
        clk), .Q(), .QN(n165) );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(AddKeyXOR1_XORInst_0_2_n1), .CK(
        clk), .Q(n203), .QN(n195) );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(AddKeyXOR1_XORInst_0_3_n1), .CK(
        clk), .Q(n216), .QN(n194) );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(AddKeyXOR1_XORInst_1_0_n1), .CK(
        clk), .Q(n204), .QN(n193) );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(AddKeyXOR1_XORInst_1_1_n1), .CK(
        clk), .Q(), .QN(n166) );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(AddKeyXOR1_XORInst_1_2_n1), .CK(
        clk), .Q(n215), .QN(n192) );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(AddKeyXOR1_XORInst_1_3_n1), .CK(
        clk), .Q(n213), .QN(n191) );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(AddKeyXOR1_XORInst_2_0_n1), .CK(
        clk), .Q(n202), .QN(n190) );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(AddKeyXOR1_XORInst_2_1_n1), .CK(
        clk), .Q(), .QN(n167) );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(AddKeyXOR1_XORInst_2_2_n1), 
        .CK(clk), .Q(n220), .QN(n189) );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(AddKeyXOR1_XORInst_2_3_n1), 
        .CK(clk), .Q(n214), .QN(n188) );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(AddKeyXOR1_XORInst_3_0_n1), 
        .CK(clk), .Q(n208), .QN(n187) );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(AddKeyXOR1_XORInst_3_1_n1), 
        .CK(clk), .Q(), .QN(n168) );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(AddKeyXOR1_XORInst_3_2_n1), 
        .CK(clk), .Q(n209), .QN(n186) );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(AddKeyXOR1_XORInst_3_3_n1), 
        .CK(clk), .Q(n201), .QN(n185) );
  DFF_X1 StateReg2_s_current_state_reg_0_ ( .D(AddKeyXOR2_XORInst_0_0_n1), 
        .CK(clk), .Q(n218), .QN(n184) );
  DFF_X1 StateReg2_s_current_state_reg_1_ ( .D(AddKeyXOR2_XORInst_0_1_n1), 
        .CK(clk), .Q(n211), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_2_ ( .D(AddKeyXOR2_XORInst_0_2_n1), 
        .CK(clk), .Q(n206), .QN(n183) );
  DFF_X1 StateReg2_s_current_state_reg_3_ ( .D(AddKeyXOR2_XORInst_0_3_n1), 
        .CK(clk), .Q(n199), .QN(n182) );
  DFF_X1 StateReg2_s_current_state_reg_4_ ( .D(AddKeyXOR2_XORInst_1_0_n1), 
        .CK(clk), .Q(n219), .QN(n181) );
  DFF_X1 StateReg2_s_current_state_reg_5_ ( .D(AddKeyXOR2_XORInst_1_1_n1), 
        .CK(clk), .Q(n212), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_6_ ( .D(AddKeyXOR2_XORInst_1_2_n1), 
        .CK(clk), .Q(n207), .QN(n180) );
  DFF_X1 StateReg2_s_current_state_reg_7_ ( .D(AddKeyXOR2_XORInst_1_3_n1), 
        .CK(clk), .Q(n200), .QN(n179) );
  DFF_X1 StateReg2_s_current_state_reg_8_ ( .D(AddKeyXOR2_XORInst_2_0_n1), 
        .CK(clk), .Q(), .QN(n178) );
  DFF_X1 StateReg2_s_current_state_reg_9_ ( .D(AddKeyXOR2_XORInst_2_1_n1), 
        .CK(clk), .Q(n221), .QN(n171) );
  DFF_X1 StateReg2_s_current_state_reg_10_ ( .D(AddKeyXOR2_XORInst_2_2_n1), 
        .CK(clk), .Q(n222), .QN(n177) );
  DFF_X1 StateReg2_s_current_state_reg_11_ ( .D(AddKeyXOR2_XORInst_2_3_n1), 
        .CK(clk), .Q(), .QN(n176) );
  DFF_X1 StateReg2_s_current_state_reg_12_ ( .D(AddKeyXOR2_XORInst_3_0_n1), 
        .CK(clk), .Q(n217), .QN(n175) );
  DFF_X1 StateReg2_s_current_state_reg_13_ ( .D(AddKeyXOR2_XORInst_3_1_n1), 
        .CK(clk), .Q(n210), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_14_ ( .D(AddKeyXOR2_XORInst_3_2_n1), 
        .CK(clk), .Q(n205), .QN(n174) );
  DFF_X1 StateReg2_s_current_state_reg_15_ ( .D(AddKeyXOR2_XORInst_3_3_n1), 
        .CK(clk), .Q(n198), .QN(n173) );
  XOR2_X1 U214 ( .A(Input[0]), .B(Key[0]), .Z(AddKeyXOR1_XORInst_0_0_n1) );
  XOR2_X1 U215 ( .A(Input[1]), .B(Key[1]), .Z(AddKeyXOR1_XORInst_0_1_n1) );
  XOR2_X1 U216 ( .A(Input[2]), .B(Key[2]), .Z(AddKeyXOR1_XORInst_0_2_n1) );
  XOR2_X1 U217 ( .A(Input[3]), .B(Key[3]), .Z(AddKeyXOR1_XORInst_0_3_n1) );
  XOR2_X1 U218 ( .A(Input[4]), .B(Key[4]), .Z(AddKeyXOR1_XORInst_1_0_n1) );
  XOR2_X1 U219 ( .A(Input[5]), .B(Key[5]), .Z(AddKeyXOR1_XORInst_1_1_n1) );
  XOR2_X1 U220 ( .A(Input[6]), .B(Key[6]), .Z(AddKeyXOR1_XORInst_1_2_n1) );
  XOR2_X1 U221 ( .A(Input[7]), .B(Key[7]), .Z(AddKeyXOR1_XORInst_1_3_n1) );
  XNOR2_X1 U222 ( .A(Input[0]), .B(Key[8]), .ZN(n223) );
  XNOR2_X1 U223 ( .A(n223), .B(Input[8]), .ZN(AddKeyXOR1_XORInst_2_0_n1) );
  XNOR2_X1 U224 ( .A(Input[1]), .B(Key[9]), .ZN(n224) );
  XNOR2_X1 U225 ( .A(n224), .B(Input[9]), .ZN(AddKeyXOR1_XORInst_2_1_n1) );
  XNOR2_X1 U226 ( .A(Input[2]), .B(Key[10]), .ZN(n225) );
  XNOR2_X1 U227 ( .A(n225), .B(Input[10]), .ZN(AddKeyXOR1_XORInst_2_2_n1) );
  XNOR2_X1 U228 ( .A(Input[3]), .B(Key[11]), .ZN(n226) );
  XNOR2_X1 U229 ( .A(n226), .B(Input[11]), .ZN(AddKeyXOR1_XORInst_2_3_n1) );
  XOR2_X1 U230 ( .A(Input[4]), .B(Input[12]), .Z(n228) );
  XNOR2_X1 U231 ( .A(Input[0]), .B(Key[12]), .ZN(n227) );
  XNOR2_X1 U232 ( .A(n228), .B(n227), .ZN(AddKeyXOR1_XORInst_3_0_n1) );
  XOR2_X1 U233 ( .A(Input[5]), .B(Input[13]), .Z(n230) );
  XNOR2_X1 U234 ( .A(Input[1]), .B(Key[13]), .ZN(n229) );
  XNOR2_X1 U235 ( .A(n230), .B(n229), .ZN(AddKeyXOR1_XORInst_3_1_n1) );
  XOR2_X1 U236 ( .A(Input[6]), .B(Input[14]), .Z(n232) );
  XNOR2_X1 U237 ( .A(Input[2]), .B(Key[14]), .ZN(n231) );
  XNOR2_X1 U238 ( .A(n232), .B(n231), .ZN(AddKeyXOR1_XORInst_3_2_n1) );
  XOR2_X1 U239 ( .A(Input[7]), .B(Input[15]), .Z(n234) );
  XNOR2_X1 U240 ( .A(Input[3]), .B(Key[15]), .ZN(n233) );
  XNOR2_X1 U241 ( .A(n234), .B(n233), .ZN(AddKeyXOR1_XORInst_3_3_n1) );
  NAND2_X1 U242 ( .A1(n216), .A2(n203), .ZN(n244) );
  NAND2_X1 U243 ( .A1(n195), .A2(n194), .ZN(n235) );
  NAND2_X1 U244 ( .A1(n235), .A2(n197), .ZN(n236) );
  NAND2_X1 U245 ( .A1(n236), .A2(n165), .ZN(n237) );
  NAND2_X1 U246 ( .A1(n244), .A2(n237), .ZN(n281) );
  XNOR2_X1 U247 ( .A(Key[16]), .B(n281), .ZN(AddKeyXOR2_XORInst_0_0_n1) );
  NAND2_X1 U248 ( .A1(n197), .A2(n203), .ZN(n240) );
  NAND2_X1 U249 ( .A1(n196), .A2(n195), .ZN(n238) );
  NAND2_X1 U250 ( .A1(n238), .A2(n194), .ZN(n239) );
  NAND2_X1 U251 ( .A1(n240), .A2(n239), .ZN(n292) );
  XOR2_X1 U252 ( .A(Key[17]), .B(n292), .Z(AddKeyXOR2_XORInst_0_1_n1) );
  NOR2_X1 U253 ( .A1(n216), .A2(n197), .ZN(n246) );
  NOR2_X1 U254 ( .A1(n194), .A2(n196), .ZN(n241) );
  NOR2_X1 U255 ( .A1(n203), .A2(n241), .ZN(n242) );
  NOR2_X1 U256 ( .A1(n165), .A2(n242), .ZN(n243) );
  NOR2_X1 U257 ( .A1(n246), .A2(n243), .ZN(n304) );
  XNOR2_X1 U258 ( .A(n304), .B(Key[18]), .ZN(AddKeyXOR2_XORInst_0_2_n1) );
  AND2_X1 U259 ( .A1(n165), .A2(n244), .ZN(n245) );
  NOR2_X1 U260 ( .A1(n246), .A2(n245), .ZN(n312) );
  XNOR2_X1 U261 ( .A(n312), .B(Key[19]), .ZN(AddKeyXOR2_XORInst_0_3_n1) );
  NOR2_X1 U262 ( .A1(n191), .A2(n192), .ZN(n259) );
  INV_X1 U263 ( .A(n259), .ZN(n250) );
  NAND2_X1 U264 ( .A1(n192), .A2(n191), .ZN(n247) );
  NAND2_X1 U265 ( .A1(n247), .A2(n204), .ZN(n248) );
  NAND2_X1 U266 ( .A1(n248), .A2(n166), .ZN(n249) );
  NAND2_X1 U267 ( .A1(n250), .A2(n249), .ZN(n287) );
  XNOR2_X1 U268 ( .A(Key[20]), .B(n287), .ZN(AddKeyXOR2_XORInst_1_0_n1) );
  NAND2_X1 U269 ( .A1(n213), .A2(n192), .ZN(n251) );
  NAND2_X1 U270 ( .A1(n251), .A2(n204), .ZN(n253) );
  NAND2_X1 U271 ( .A1(n215), .A2(n191), .ZN(n252) );
  NAND2_X1 U272 ( .A1(n253), .A2(n252), .ZN(n296) );
  XOR2_X1 U273 ( .A(n296), .B(Key[21]), .Z(AddKeyXOR2_XORInst_1_1_n1) );
  NOR2_X1 U274 ( .A1(n213), .A2(n204), .ZN(n257) );
  NOR2_X1 U275 ( .A1(n191), .A2(n193), .ZN(n254) );
  NOR2_X1 U276 ( .A1(n215), .A2(n254), .ZN(n255) );
  NOR2_X1 U277 ( .A1(n166), .A2(n255), .ZN(n256) );
  NOR2_X1 U278 ( .A1(n257), .A2(n256), .ZN(n297) );
  XNOR2_X1 U279 ( .A(n297), .B(Key[22]), .ZN(AddKeyXOR2_XORInst_1_2_n1) );
  NOR2_X1 U280 ( .A1(n166), .A2(n257), .ZN(n258) );
  NOR2_X1 U281 ( .A1(n259), .A2(n258), .ZN(n305) );
  XOR2_X1 U282 ( .A(n305), .B(Key[23]), .Z(AddKeyXOR2_XORInst_1_3_n1) );
  NAND2_X1 U283 ( .A1(n189), .A2(n188), .ZN(n260) );
  NAND2_X1 U284 ( .A1(n260), .A2(n202), .ZN(n261) );
  NAND2_X1 U285 ( .A1(n261), .A2(n167), .ZN(n263) );
  NOR2_X1 U286 ( .A1(n188), .A2(n189), .ZN(n278) );
  INV_X1 U287 ( .A(n278), .ZN(n262) );
  NAND2_X1 U288 ( .A1(n263), .A2(n262), .ZN(n264) );
  XNOR2_X1 U289 ( .A(n264), .B(n281), .ZN(n265) );
  XNOR2_X1 U290 ( .A(Key[24]), .B(n265), .ZN(AddKeyXOR2_XORInst_2_0_n1) );
  NAND2_X1 U291 ( .A1(n214), .A2(n190), .ZN(n266) );
  NAND2_X1 U292 ( .A1(n266), .A2(n220), .ZN(n268) );
  NAND2_X1 U293 ( .A1(n202), .A2(n188), .ZN(n267) );
  NAND2_X1 U294 ( .A1(n268), .A2(n267), .ZN(n269) );
  XNOR2_X1 U295 ( .A(n269), .B(n292), .ZN(n270) );
  XNOR2_X1 U296 ( .A(Key[25]), .B(n270), .ZN(AddKeyXOR2_XORInst_2_1_n1) );
  XNOR2_X1 U297 ( .A(Key[26]), .B(n304), .ZN(n275) );
  NOR2_X1 U298 ( .A1(n214), .A2(n202), .ZN(n276) );
  NOR2_X1 U299 ( .A1(n188), .A2(n190), .ZN(n271) );
  NOR2_X1 U300 ( .A1(n220), .A2(n271), .ZN(n272) );
  NOR2_X1 U301 ( .A1(n167), .A2(n272), .ZN(n273) );
  NOR2_X1 U302 ( .A1(n276), .A2(n273), .ZN(n274) );
  XNOR2_X1 U303 ( .A(n275), .B(n274), .ZN(AddKeyXOR2_XORInst_2_2_n1) );
  NOR2_X1 U304 ( .A1(n167), .A2(n276), .ZN(n277) );
  NOR2_X1 U305 ( .A1(n278), .A2(n277), .ZN(n279) );
  XOR2_X1 U306 ( .A(n312), .B(n279), .Z(n280) );
  XNOR2_X1 U307 ( .A(Key[27]), .B(n280), .ZN(AddKeyXOR2_XORInst_2_3_n1) );
  XNOR2_X1 U308 ( .A(n281), .B(Key[28]), .ZN(n286) );
  NAND2_X1 U309 ( .A1(n201), .A2(n209), .ZN(n307) );
  NAND2_X1 U310 ( .A1(n186), .A2(n185), .ZN(n282) );
  NAND2_X1 U311 ( .A1(n282), .A2(n208), .ZN(n283) );
  NAND2_X1 U312 ( .A1(n283), .A2(n168), .ZN(n284) );
  NAND2_X1 U313 ( .A1(n307), .A2(n284), .ZN(n285) );
  XNOR2_X1 U314 ( .A(n286), .B(n285), .ZN(n288) );
  XNOR2_X1 U315 ( .A(n288), .B(n287), .ZN(AddKeyXOR2_XORInst_3_0_n1) );
  NAND2_X1 U316 ( .A1(n201), .A2(n187), .ZN(n289) );
  NAND2_X1 U317 ( .A1(n289), .A2(n209), .ZN(n291) );
  NAND2_X1 U318 ( .A1(n208), .A2(n185), .ZN(n290) );
  NAND2_X1 U319 ( .A1(n291), .A2(n290), .ZN(n293) );
  XNOR2_X1 U320 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U321 ( .A(Key[29]), .B(n294), .Z(n295) );
  XNOR2_X1 U322 ( .A(n296), .B(n295), .ZN(AddKeyXOR2_XORInst_3_1_n1) );
  XNOR2_X1 U323 ( .A(n297), .B(Key[30]), .ZN(n302) );
  NOR2_X1 U324 ( .A1(n201), .A2(n208), .ZN(n306) );
  NOR2_X1 U325 ( .A1(n185), .A2(n187), .ZN(n298) );
  NOR2_X1 U326 ( .A1(n209), .A2(n298), .ZN(n299) );
  NOR2_X1 U327 ( .A1(n168), .A2(n299), .ZN(n300) );
  NOR2_X1 U328 ( .A1(n306), .A2(n300), .ZN(n301) );
  XNOR2_X1 U329 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U330 ( .A(n304), .B(n303), .ZN(AddKeyXOR2_XORInst_3_2_n1) );
  XOR2_X1 U331 ( .A(Key[31]), .B(n305), .Z(n310) );
  OR2_X1 U332 ( .A1(n168), .A2(n306), .ZN(n308) );
  NAND2_X1 U333 ( .A1(n308), .A2(n307), .ZN(n309) );
  XNOR2_X1 U334 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U335 ( .A(n312), .B(n311), .ZN(AddKeyXOR2_XORInst_3_3_n1) );
  NOR2_X1 U336 ( .A1(n182), .A2(n183), .ZN(n339) );
  NOR2_X1 U337 ( .A1(n206), .A2(n199), .ZN(n313) );
  NOR2_X1 U338 ( .A1(n184), .A2(n313), .ZN(n314) );
  NOR2_X1 U339 ( .A1(n314), .A2(n211), .ZN(n315) );
  NOR2_X1 U340 ( .A1(n339), .A2(n315), .ZN(Output[0]) );
  NAND2_X1 U341 ( .A1(n178), .A2(n176), .ZN(n320) );
  NOR2_X1 U342 ( .A1(n178), .A2(n176), .ZN(n316) );
  NOR2_X1 U343 ( .A1(n222), .A2(n316), .ZN(n317) );
  OR2_X1 U344 ( .A1(n171), .A2(n317), .ZN(n318) );
  NAND2_X1 U345 ( .A1(n320), .A2(n318), .ZN(Output[10]) );
  NOR2_X1 U346 ( .A1(n176), .A2(n177), .ZN(n356) );
  OR2_X1 U347 ( .A1(n356), .A2(n221), .ZN(n319) );
  NAND2_X1 U348 ( .A1(n320), .A2(n319), .ZN(Output[11]) );
  NOR2_X1 U349 ( .A1(n173), .A2(n174), .ZN(n330) );
  NOR2_X1 U350 ( .A1(n205), .A2(n198), .ZN(n321) );
  NOR2_X1 U351 ( .A1(n175), .A2(n321), .ZN(n322) );
  NOR2_X1 U352 ( .A1(n322), .A2(n210), .ZN(n323) );
  NOR2_X1 U353 ( .A1(n330), .A2(n323), .ZN(Output[12]) );
  NAND2_X1 U354 ( .A1(n217), .A2(n205), .ZN(n326) );
  NAND2_X1 U355 ( .A1(n175), .A2(n174), .ZN(n324) );
  NAND2_X1 U356 ( .A1(n324), .A2(n173), .ZN(n325) );
  NAND2_X1 U357 ( .A1(n326), .A2(n325), .ZN(Output[13]) );
  NAND2_X1 U358 ( .A1(n173), .A2(n175), .ZN(n332) );
  NAND2_X1 U359 ( .A1(n217), .A2(n198), .ZN(n327) );
  NAND2_X1 U360 ( .A1(n327), .A2(n174), .ZN(n328) );
  NAND2_X1 U361 ( .A1(n328), .A2(n210), .ZN(n329) );
  NAND2_X1 U362 ( .A1(n332), .A2(n329), .ZN(Output[14]) );
  OR2_X1 U363 ( .A1(n330), .A2(n210), .ZN(n331) );
  NAND2_X1 U364 ( .A1(n332), .A2(n331), .ZN(Output[15]) );
  NAND2_X1 U365 ( .A1(n218), .A2(n206), .ZN(n335) );
  NAND2_X1 U366 ( .A1(n184), .A2(n183), .ZN(n333) );
  NAND2_X1 U367 ( .A1(n333), .A2(n182), .ZN(n334) );
  NAND2_X1 U368 ( .A1(n335), .A2(n334), .ZN(Output[1]) );
  NAND2_X1 U369 ( .A1(n182), .A2(n184), .ZN(n341) );
  NAND2_X1 U370 ( .A1(n218), .A2(n199), .ZN(n336) );
  NAND2_X1 U371 ( .A1(n336), .A2(n183), .ZN(n337) );
  NAND2_X1 U372 ( .A1(n337), .A2(n211), .ZN(n338) );
  NAND2_X1 U373 ( .A1(n341), .A2(n338), .ZN(Output[2]) );
  OR2_X1 U374 ( .A1(n339), .A2(n211), .ZN(n340) );
  NAND2_X1 U375 ( .A1(n341), .A2(n340), .ZN(Output[3]) );
  NOR2_X1 U376 ( .A1(n179), .A2(n180), .ZN(n351) );
  NOR2_X1 U377 ( .A1(n207), .A2(n200), .ZN(n342) );
  NOR2_X1 U378 ( .A1(n181), .A2(n342), .ZN(n343) );
  NOR2_X1 U379 ( .A1(n343), .A2(n212), .ZN(n344) );
  NOR2_X1 U380 ( .A1(n351), .A2(n344), .ZN(Output[4]) );
  NAND2_X1 U381 ( .A1(n219), .A2(n207), .ZN(n347) );
  NAND2_X1 U382 ( .A1(n181), .A2(n180), .ZN(n345) );
  NAND2_X1 U383 ( .A1(n345), .A2(n179), .ZN(n346) );
  NAND2_X1 U384 ( .A1(n347), .A2(n346), .ZN(Output[5]) );
  NAND2_X1 U385 ( .A1(n179), .A2(n181), .ZN(n353) );
  NAND2_X1 U386 ( .A1(n219), .A2(n200), .ZN(n348) );
  NAND2_X1 U387 ( .A1(n348), .A2(n180), .ZN(n349) );
  NAND2_X1 U388 ( .A1(n349), .A2(n212), .ZN(n350) );
  NAND2_X1 U389 ( .A1(n353), .A2(n350), .ZN(Output[6]) );
  OR2_X1 U390 ( .A1(n351), .A2(n212), .ZN(n352) );
  NAND2_X1 U391 ( .A1(n353), .A2(n352), .ZN(Output[7]) );
  AND2_X1 U392 ( .A1(n176), .A2(n177), .ZN(n354) );
  NOR2_X1 U393 ( .A1(n178), .A2(n354), .ZN(n355) );
  NOR2_X1 U394 ( .A1(n221), .A2(n355), .ZN(n357) );
  NOR2_X1 U395 ( .A1(n357), .A2(n356), .ZN(Output[8]) );
  OR2_X1 U396 ( .A1(n177), .A2(n178), .ZN(n360) );
  NAND2_X1 U397 ( .A1(n177), .A2(n178), .ZN(n358) );
  NAND2_X1 U398 ( .A1(n358), .A2(n176), .ZN(n359) );
  NAND2_X1 U399 ( .A1(n360), .A2(n359), .ZN(Output[9]) );
endmodule

