
module Cipher ( clk, rst, EncDec, Input, Key, Output );
  input [63:0] Input;
  input [63:0] Key;
  output [63:0] Output;
  (* fiver="clock" *)input clk;
  (* fiver="control" *)input rst;
  (* fiver="control" *)input EncDec;
  wire   MCOutput_63_, MCOutput_62_, MCOutput_61_, MCOutput_60_, MCOutput_59_,
         MCOutput_58_, MCOutput_57_, MCOutput_56_, MCOutput_55_, MCOutput_54_,
         MCOutput_53_, MCOutput_52_, MCOutput_51_, MCOutput_50_, MCOutput_49_,
         MCOutput_48_, MCOutput_47_, MCOutput_46_, MCOutput_45_, MCOutput_44_,
         MCOutput_43_, MCOutput_42_, MCOutput_41_, MCOutput_40_, MCOutput_39_,
         MCOutput_38_, MCOutput_37_, MCOutput_36_, MCOutput_35_, MCOutput_34_,
         MCOutput_33_, MCOutput_32_, MCInst_XOR_r0_Inst_0_n5,
         MCInst_XOR_r0_Inst_1_n5, MCInst_XOR_r0_Inst_2_n5,
         MCInst_XOR_r0_Inst_3_n5, MCInst_XOR_r0_Inst_4_n5,
         MCInst_XOR_r0_Inst_5_n5, MCInst_XOR_r0_Inst_6_n5,
         MCInst_XOR_r0_Inst_7_n5, MCInst_XOR_r0_Inst_8_n5,
         MCInst_XOR_r0_Inst_9_n5, MCInst_XOR_r0_Inst_10_n5,
         MCInst_XOR_r0_Inst_11_n5, MCInst_XOR_r0_Inst_12_n5,
         MCInst_XOR_r0_Inst_13_n5, MCInst_XOR_r0_Inst_14_n5,
         MCInst_XOR_r0_Inst_15_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n17,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n18,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n38,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n37,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n16,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n15,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n14,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n13,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n12,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n11,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n10,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n9,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n8,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n7,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n6,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n5,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n4,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n3,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n2,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n1,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n35,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n34,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n33,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n32,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n31,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n30,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n29,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n28,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n27,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n26,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n25,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n24,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n23,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n22,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n21,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n20,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n19,
         SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n18,
         Red_PlaintextInst_LFInst_0_LFInst_0_n3,
         Red_PlaintextInst_LFInst_0_LFInst_1_n3,
         Red_PlaintextInst_LFInst_0_LFInst_2_n3,
         Red_PlaintextInst_LFInst_1_LFInst_0_n3,
         Red_PlaintextInst_LFInst_1_LFInst_1_n3,
         Red_PlaintextInst_LFInst_1_LFInst_2_n3,
         Red_PlaintextInst_LFInst_2_LFInst_0_n3,
         Red_PlaintextInst_LFInst_2_LFInst_1_n3,
         Red_PlaintextInst_LFInst_2_LFInst_2_n3,
         Red_PlaintextInst_LFInst_3_LFInst_0_n3,
         Red_PlaintextInst_LFInst_3_LFInst_1_n3,
         Red_PlaintextInst_LFInst_3_LFInst_2_n3,
         Red_PlaintextInst_LFInst_4_LFInst_0_n3,
         Red_PlaintextInst_LFInst_4_LFInst_1_n3,
         Red_PlaintextInst_LFInst_4_LFInst_2_n3,
         Red_PlaintextInst_LFInst_5_LFInst_0_n3,
         Red_PlaintextInst_LFInst_5_LFInst_1_n3,
         Red_PlaintextInst_LFInst_5_LFInst_2_n3,
         Red_PlaintextInst_LFInst_6_LFInst_0_n3,
         Red_PlaintextInst_LFInst_6_LFInst_1_n3,
         Red_PlaintextInst_LFInst_6_LFInst_2_n3,
         Red_PlaintextInst_LFInst_7_LFInst_0_n3,
         Red_PlaintextInst_LFInst_7_LFInst_1_n3,
         Red_PlaintextInst_LFInst_7_LFInst_2_n3,
         Red_PlaintextInst_LFInst_8_LFInst_0_n3,
         Red_PlaintextInst_LFInst_8_LFInst_1_n3,
         Red_PlaintextInst_LFInst_8_LFInst_2_n3,
         Red_PlaintextInst_LFInst_9_LFInst_0_n3,
         Red_PlaintextInst_LFInst_9_LFInst_1_n3,
         Red_PlaintextInst_LFInst_9_LFInst_2_n3,
         Red_PlaintextInst_LFInst_10_LFInst_0_n3,
         Red_PlaintextInst_LFInst_10_LFInst_1_n3,
         Red_PlaintextInst_LFInst_10_LFInst_2_n3,
         Red_PlaintextInst_LFInst_11_LFInst_0_n3,
         Red_PlaintextInst_LFInst_11_LFInst_1_n3,
         Red_PlaintextInst_LFInst_11_LFInst_2_n3,
         Red_PlaintextInst_LFInst_12_LFInst_0_n3,
         Red_PlaintextInst_LFInst_12_LFInst_1_n3,
         Red_PlaintextInst_LFInst_12_LFInst_2_n3,
         Red_PlaintextInst_LFInst_13_LFInst_0_n3,
         Red_PlaintextInst_LFInst_13_LFInst_1_n3,
         Red_PlaintextInst_LFInst_13_LFInst_2_n3,
         Red_PlaintextInst_LFInst_14_LFInst_0_n3,
         Red_PlaintextInst_LFInst_14_LFInst_1_n3,
         Red_PlaintextInst_LFInst_14_LFInst_2_n3,
         Red_PlaintextInst_LFInst_15_LFInst_0_n3,
         Red_PlaintextInst_LFInst_15_LFInst_1_n3,
         Red_PlaintextInst_LFInst_15_LFInst_2_n3, Red_MCInst_XOR_r0_Inst_0_n5,
         Red_MCInst_XOR_r0_Inst_1_n5, Red_MCInst_XOR_r0_Inst_2_n5,
         Red_MCInst_XOR_r0_Inst_3_n5, Red_MCInst_XOR_r0_Inst_4_n5,
         Red_MCInst_XOR_r0_Inst_5_n5, Red_MCInst_XOR_r0_Inst_6_n5,
         Red_MCInst_XOR_r0_Inst_7_n5, Red_MCInst_XOR_r0_Inst_8_n5,
         Red_MCInst_XOR_r0_Inst_9_n5, Red_MCInst_XOR_r0_Inst_10_n5,
         Red_MCInst_XOR_r0_Inst_11_n5,
         StateRegOutputF_inst_LFInst_0_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_0_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_0_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_1_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_1_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_1_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_2_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_2_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_2_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_3_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_3_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_3_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_4_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_4_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_4_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_5_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_5_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_5_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_6_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_6_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_6_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_7_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_7_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_7_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_8_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_8_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_8_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_9_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_9_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_9_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_10_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_10_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_10_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_11_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_11_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_11_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_12_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_12_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_12_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_13_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_13_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_13_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_14_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_14_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_14_LFInst_2_n3,
         StateRegOutputF_inst_LFInst_15_LFInst_0_n3,
         StateRegOutputF_inst_LFInst_15_LFInst_1_n3,
         StateRegOutputF_inst_LFInst_15_LFInst_2_n3,
         CipherErrorVecGen_XORInst_0_0_n6, CipherErrorVecGen_XORInst_0_1_n5,
         CipherErrorVecGen_XORInst_0_2_n2, CipherErrorVecGen_XORInst_1_0_n6,
         CipherErrorVecGen_XORInst_1_1_n5, CipherErrorVecGen_XORInst_1_2_n2,
         CipherErrorVecGen_XORInst_2_0_n6, CipherErrorVecGen_XORInst_2_1_n5,
         CipherErrorVecGen_XORInst_2_2_n2, CipherErrorVecGen_XORInst_3_0_n6,
         CipherErrorVecGen_XORInst_3_1_n2, CipherErrorVecGen_XORInst_3_2_n2,
         CipherErrorVecGen_XORInst_4_0_n6, CipherErrorVecGen_XORInst_4_1_n5,
         CipherErrorVecGen_XORInst_4_2_n2, CipherErrorVecGen_XORInst_5_0_n6,
         CipherErrorVecGen_XORInst_5_1_n5, CipherErrorVecGen_XORInst_5_2_n2,
         CipherErrorVecGen_XORInst_6_0_n6, CipherErrorVecGen_XORInst_6_1_n5,
         CipherErrorVecGen_XORInst_6_2_n2, CipherErrorVecGen_XORInst_7_0_n6,
         CipherErrorVecGen_XORInst_7_1_n5, CipherErrorVecGen_XORInst_7_2_n2,
         CipherErrorVecGen_XORInst_8_0_n6, CipherErrorVecGen_XORInst_8_1_n5,
         CipherErrorVecGen_XORInst_8_2_n2, CipherErrorVecGen_XORInst_9_0_n6,
         CipherErrorVecGen_XORInst_9_1_n5, CipherErrorVecGen_XORInst_9_2_n2,
         CipherErrorVecGen_XORInst_10_0_n6, CipherErrorVecGen_XORInst_10_1_n5,
         CipherErrorVecGen_XORInst_10_2_n2, CipherErrorVecGen_XORInst_11_0_n6,
         CipherErrorVecGen_XORInst_11_1_n5, CipherErrorVecGen_XORInst_11_2_n2,
         CipherErrorVecGen_XORInst_12_0_n6, CipherErrorVecGen_XORInst_12_1_n5,
         CipherErrorVecGen_XORInst_12_2_n2, CipherErrorVecGen_XORInst_13_0_n6,
         CipherErrorVecGen_XORInst_13_1_n5, CipherErrorVecGen_XORInst_13_2_n2,
         CipherErrorVecGen_XORInst_14_0_n6, CipherErrorVecGen_XORInst_14_1_n5,
         CipherErrorVecGen_XORInst_14_2_n2, CipherErrorVecGen_XORInst_15_0_n6,
         CipherErrorVecGen_XORInst_15_1_n5, CipherErrorVecGen_XORInst_15_2_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n1,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n2,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n19,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n18,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n17,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n16,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n15,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n14,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n13,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n12,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n11,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n10,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n9,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n8,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n7,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n6,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n5,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n4,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n3,
         SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n2,
         StateRegOutputF_inst2_LFInst_0_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_0_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_0_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_1_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_1_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_1_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_2_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_2_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_2_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_3_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_3_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_3_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_4_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_4_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_4_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_5_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_5_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_5_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_6_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_6_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_6_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_7_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_7_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_7_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_8_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_8_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_8_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_9_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_9_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_9_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_10_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_10_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_10_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_11_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_11_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_11_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_12_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_12_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_12_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_13_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_13_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_13_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_14_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_14_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_14_LFInst_2_n3,
         StateRegOutputF_inst2_LFInst_15_LFInst_0_n3,
         StateRegOutputF_inst2_LFInst_15_LFInst_1_n3,
         StateRegOutputF_inst2_LFInst_15_LFInst_2_n3,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n39,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n46,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n45,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n44,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n43,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n42,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n41,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n40,
         SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n39,
         Red_K1Inst_LFInst_0_LFInst_0_n3, Red_K1Inst_LFInst_0_LFInst_1_n3,
         Red_K1Inst_LFInst_0_LFInst_2_n3, Red_K1Inst_LFInst_1_LFInst_0_n3,
         Red_K1Inst_LFInst_1_LFInst_1_n3, Red_K1Inst_LFInst_1_LFInst_2_n3,
         Red_K1Inst_LFInst_2_LFInst_0_n3, Red_K1Inst_LFInst_2_LFInst_1_n3,
         Red_K1Inst_LFInst_2_LFInst_2_n3, Red_K1Inst_LFInst_3_LFInst_0_n3,
         Red_K1Inst_LFInst_3_LFInst_1_n3, Red_K1Inst_LFInst_3_LFInst_2_n3,
         Red_K1Inst_LFInst_4_LFInst_0_n3, Red_K1Inst_LFInst_4_LFInst_1_n3,
         Red_K1Inst_LFInst_4_LFInst_2_n3, Red_K1Inst_LFInst_5_LFInst_0_n3,
         Red_K1Inst_LFInst_5_LFInst_1_n3, Red_K1Inst_LFInst_5_LFInst_2_n3,
         Red_K1Inst_LFInst_6_LFInst_0_n3, Red_K1Inst_LFInst_6_LFInst_1_n3,
         Red_K1Inst_LFInst_6_LFInst_2_n3, Red_K1Inst_LFInst_7_LFInst_0_n3,
         Red_K1Inst_LFInst_7_LFInst_1_n3, Red_K1Inst_LFInst_7_LFInst_2_n3,
         Red_K1Inst_LFInst_8_LFInst_0_n3, Red_K1Inst_LFInst_8_LFInst_1_n3,
         Red_K1Inst_LFInst_8_LFInst_2_n3, Red_K1Inst_LFInst_9_LFInst_0_n3,
         Red_K1Inst_LFInst_9_LFInst_1_n3, Red_K1Inst_LFInst_9_LFInst_2_n3,
         Red_K1Inst_LFInst_10_LFInst_0_n3, Red_K1Inst_LFInst_10_LFInst_1_n3,
         Red_K1Inst_LFInst_10_LFInst_2_n3, Red_K1Inst_LFInst_11_LFInst_0_n3,
         Red_K1Inst_LFInst_11_LFInst_1_n3, Red_K1Inst_LFInst_11_LFInst_2_n3,
         Red_K1Inst_LFInst_12_LFInst_0_n3, Red_K1Inst_LFInst_12_LFInst_1_n3,
         Red_K1Inst_LFInst_12_LFInst_2_n3, Red_K1Inst_LFInst_13_LFInst_0_n3,
         Red_K1Inst_LFInst_13_LFInst_1_n3, Red_K1Inst_LFInst_13_LFInst_2_n3,
         Red_K1Inst_LFInst_14_LFInst_0_n3, Red_K1Inst_LFInst_14_LFInst_1_n3,
         Red_K1Inst_LFInst_14_LFInst_2_n3, Red_K1Inst_LFInst_15_LFInst_0_n3,
         Red_K1Inst_LFInst_15_LFInst_1_n3, Red_K1Inst_LFInst_15_LFInst_2_n3;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] StateRegOutput;
  wire   [47:0] CipherErrorVec;
  wire   [63:0] Feedback;
  wire   [47:24] Red_Input;
  wire   [47:0] Red_MCOutput;
  wire   [47:0] Red_AddRoundKeyOutput;
  wire   [47:0] Red_K1;
  wire   [47:0] Red_StateRegOutput;
  wire   [47:0] StateRegOutputF;
  wire   [47:0] Red_Feedback;
  wire   [47:0] FeedbackF;
  wire   [47:0] CipherErrorVec2;

  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2 ( .A(MCInst_XOR_r0_Inst_0_n5), .B(Input[16]), .ZN(MCOutput_48_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U1 ( .A(Input[0]), .B(Input[48]), .ZN(
        MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_0_U1 ( .A(Input[32]), .B(Input[0]), .Z(
        MCOutput_32_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2 ( .A(MCInst_XOR_r0_Inst_1_n5), .B(Input[17]), .ZN(MCOutput_49_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U1 ( .A(Input[1]), .B(Input[49]), .ZN(
        MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_1_U1 ( .A(Input[33]), .B(Input[1]), .Z(
        MCOutput_33_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2 ( .A(MCInst_XOR_r0_Inst_2_n5), .B(Input[18]), .ZN(MCOutput_50_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U1 ( .A(Input[2]), .B(Input[50]), .ZN(
        MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_2_U1 ( .A(Input[34]), .B(Input[2]), .Z(
        MCOutput_34_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2 ( .A(MCInst_XOR_r0_Inst_3_n5), .B(Input[19]), .ZN(MCOutput_51_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U1 ( .A(Input[3]), .B(Input[51]), .ZN(
        MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_3_U1 ( .A(Input[35]), .B(Input[3]), .Z(
        MCOutput_35_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2 ( .A(MCInst_XOR_r0_Inst_4_n5), .B(Input[20]), .ZN(MCOutput_52_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U1 ( .A(Input[4]), .B(Input[52]), .ZN(
        MCInst_XOR_r0_Inst_4_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_4_U1 ( .A(Input[36]), .B(Input[4]), .Z(
        MCOutput_36_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2 ( .A(MCInst_XOR_r0_Inst_5_n5), .B(Input[21]), .ZN(MCOutput_53_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U1 ( .A(Input[5]), .B(Input[53]), .ZN(
        MCInst_XOR_r0_Inst_5_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_5_U1 ( .A(Input[37]), .B(Input[5]), .Z(
        MCOutput_37_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2 ( .A(MCInst_XOR_r0_Inst_6_n5), .B(Input[22]), .ZN(MCOutput_54_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U1 ( .A(Input[6]), .B(Input[54]), .ZN(
        MCInst_XOR_r0_Inst_6_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_6_U1 ( .A(Input[38]), .B(Input[6]), .Z(
        MCOutput_38_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2 ( .A(MCInst_XOR_r0_Inst_7_n5), .B(Input[23]), .ZN(MCOutput_55_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U1 ( .A(Input[7]), .B(Input[55]), .ZN(
        MCInst_XOR_r0_Inst_7_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_7_U1 ( .A(Input[39]), .B(Input[7]), .Z(
        MCOutput_39_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2 ( .A(MCInst_XOR_r0_Inst_8_n5), .B(Input[24]), .ZN(MCOutput_56_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U1 ( .A(Input[8]), .B(Input[56]), .ZN(
        MCInst_XOR_r0_Inst_8_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_8_U1 ( .A(Input[40]), .B(Input[8]), .Z(
        MCOutput_40_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2 ( .A(MCInst_XOR_r0_Inst_9_n5), .B(Input[25]), .ZN(MCOutput_57_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U1 ( .A(Input[9]), .B(Input[57]), .ZN(
        MCInst_XOR_r0_Inst_9_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_9_U1 ( .A(Input[41]), .B(Input[9]), .Z(
        MCOutput_41_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2 ( .A(MCInst_XOR_r0_Inst_10_n5), .B(
        Input[26]), .ZN(MCOutput_58_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U1 ( .A(Input[10]), .B(Input[58]), .ZN(
        MCInst_XOR_r0_Inst_10_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_10_U1 ( .A(Input[42]), .B(Input[10]), .Z(
        MCOutput_42_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2 ( .A(MCInst_XOR_r0_Inst_11_n5), .B(
        Input[27]), .ZN(MCOutput_59_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U1 ( .A(Input[11]), .B(Input[59]), .ZN(
        MCInst_XOR_r0_Inst_11_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_11_U1 ( .A(Input[43]), .B(Input[11]), .Z(
        MCOutput_43_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2 ( .A(MCInst_XOR_r0_Inst_12_n5), .B(
        Input[28]), .ZN(MCOutput_60_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U1 ( .A(Input[12]), .B(Input[60]), .ZN(
        MCInst_XOR_r0_Inst_12_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_12_U1 ( .A(Input[44]), .B(Input[12]), .Z(
        MCOutput_44_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2 ( .A(MCInst_XOR_r0_Inst_13_n5), .B(
        Input[29]), .ZN(MCOutput_61_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U1 ( .A(Input[13]), .B(Input[61]), .ZN(
        MCInst_XOR_r0_Inst_13_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_13_U1 ( .A(Input[45]), .B(Input[13]), .Z(
        MCOutput_45_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2 ( .A(MCInst_XOR_r0_Inst_14_n5), .B(
        Input[30]), .ZN(MCOutput_62_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U1 ( .A(Input[14]), .B(Input[62]), .ZN(
        MCInst_XOR_r0_Inst_14_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_14_U1 ( .A(Input[46]), .B(Input[14]), .Z(
        MCOutput_46_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2 ( .A(MCInst_XOR_r0_Inst_15_n5), .B(
        Input[31]), .ZN(MCOutput_63_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U1 ( .A(Input[15]), .B(Input[63]), .ZN(
        MCInst_XOR_r0_Inst_15_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_15_U1 ( .A(Input[47]), .B(Input[15]), .Z(
        MCOutput_47_) );
  XOR2_X1 AddKeyXOR1_XORInst_0_0_U1 ( .A(MCOutput_48_), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_1_U1 ( .A(MCOutput_49_), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_2_U1 ( .A(MCOutput_50_), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_3_U1 ( .A(MCOutput_51_), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_0_U1 ( .A(MCOutput_52_), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_1_U1 ( .A(MCOutput_53_), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_2_U1 ( .A(MCOutput_54_), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_3_U1 ( .A(MCOutput_55_), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_0_U1 ( .A(MCOutput_56_), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_1_U1 ( .A(MCOutput_57_), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_2_U1 ( .A(MCOutput_58_), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_3_U1 ( .A(MCOutput_59_), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_0_U1 ( .A(MCOutput_60_), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_1_U1 ( .A(MCOutput_61_), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_2_U1 ( .A(MCOutput_62_), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_3_U1 ( .A(MCOutput_63_), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_0_U1 ( .A(MCOutput_40_), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_1_U1 ( .A(MCOutput_41_), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_2_U1 ( .A(MCOutput_42_), .B(Key[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1 ( .A(MCOutput_43_), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_0_U1 ( .A(MCOutput_44_), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_1_U1 ( .A(MCOutput_45_), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_2_U1 ( .A(MCOutput_46_), .B(Key[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_3_U1 ( .A(MCOutput_47_), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_0_U1 ( .A(Input[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_1_U1 ( .A(Input[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_2_U1 ( .A(Input[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_3_U1 ( .A(Input[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_0_U1 ( .A(Input[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_1_U1 ( .A(Input[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_2_U1 ( .A(Input[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_3_U1 ( .A(Input[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_0_U1 ( .A(Input[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_1_U1 ( .A(Input[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_2_U1 ( .A(Input[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_3_U1 ( .A(Input[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_0_U1 ( .A(Input[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_1_U1 ( .A(Input[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_2_U1 ( .A(Input[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_3_U1 ( .A(Input[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_0_U1 ( .A(Input[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_1_U1 ( .A(Input[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_2_U1 ( .A(Input[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_3_U1 ( .A(Input[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_0_U1 ( .A(Input[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_1_U1 ( .A(Input[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_2_U1 ( .A(Input[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_3_U1 ( .A(Input[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_0_U1 ( .A(Input[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_1_U1 ( .A(Input[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_2_U1 ( .A(Input[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_3_U1 ( .A(Input[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_0_U1 ( .A(Input[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_1_U1 ( .A(Input[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_2_U1 ( .A(Input[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_3_U1 ( .A(Input[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_0_U1 ( .A(MCOutput_32_), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_1_U1 ( .A(MCOutput_33_), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_2_U1 ( .A(MCOutput_34_), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_3_U1 ( .A(MCOutput_35_), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_0_U1 ( .A(MCOutput_36_), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_1_U1 ( .A(MCOutput_37_), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_2_U1 ( .A(MCOutput_38_), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_3_U1 ( .A(MCOutput_39_), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(AddRoundKeyOutput[0]), .CK(clk), 
        .Q(StateRegOutput[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(AddRoundKeyOutput[1]), .CK(clk), 
        .Q(StateRegOutput[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(AddRoundKeyOutput[2]), .CK(clk), 
        .Q(StateRegOutput[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(AddRoundKeyOutput[3]), .CK(clk), 
        .Q(StateRegOutput[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(AddRoundKeyOutput[4]), .CK(clk), 
        .Q(StateRegOutput[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(AddRoundKeyOutput[5]), .CK(clk), 
        .Q(StateRegOutput[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(AddRoundKeyOutput[6]), .CK(clk), 
        .Q(StateRegOutput[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(AddRoundKeyOutput[7]), .CK(clk), 
        .Q(StateRegOutput[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(AddRoundKeyOutput[8]), .CK(clk), 
        .Q(StateRegOutput[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(AddRoundKeyOutput[9]), .CK(clk), 
        .Q(StateRegOutput[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(AddRoundKeyOutput[10]), .CK(clk), .Q(StateRegOutput[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(AddRoundKeyOutput[11]), .CK(clk), .Q(StateRegOutput[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(AddRoundKeyOutput[12]), .CK(clk), .Q(StateRegOutput[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(AddRoundKeyOutput[13]), .CK(clk), .Q(StateRegOutput[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(AddRoundKeyOutput[14]), .CK(clk), .Q(StateRegOutput[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(AddRoundKeyOutput[15]), .CK(clk), .Q(StateRegOutput[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(AddRoundKeyOutput[16]), .CK(clk), .Q(StateRegOutput[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(AddRoundKeyOutput[17]), .CK(clk), .Q(StateRegOutput[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(AddRoundKeyOutput[18]), .CK(clk), .Q(StateRegOutput[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(AddRoundKeyOutput[19]), .CK(clk), .Q(StateRegOutput[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(AddRoundKeyOutput[20]), .CK(clk), .Q(StateRegOutput[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(AddRoundKeyOutput[21]), .CK(clk), .Q(StateRegOutput[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(AddRoundKeyOutput[22]), .CK(clk), .Q(StateRegOutput[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(AddRoundKeyOutput[23]), .CK(clk), .Q(StateRegOutput[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(AddRoundKeyOutput[24]), .CK(clk), .Q(StateRegOutput[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(AddRoundKeyOutput[25]), .CK(clk), .Q(StateRegOutput[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(AddRoundKeyOutput[26]), .CK(clk), .Q(StateRegOutput[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(AddRoundKeyOutput[27]), .CK(clk), .Q(StateRegOutput[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(AddRoundKeyOutput[28]), .CK(clk), .Q(StateRegOutput[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(AddRoundKeyOutput[29]), .CK(clk), .Q(StateRegOutput[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(AddRoundKeyOutput[30]), .CK(clk), .Q(StateRegOutput[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(AddRoundKeyOutput[31]), .CK(clk), .Q(StateRegOutput[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(AddRoundKeyOutput[32]), .CK(clk), .Q(StateRegOutput[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(AddRoundKeyOutput[33]), .CK(clk), .Q(StateRegOutput[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(AddRoundKeyOutput[34]), .CK(clk), .Q(StateRegOutput[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(AddRoundKeyOutput[35]), .CK(clk), .Q(StateRegOutput[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(AddRoundKeyOutput[36]), .CK(clk), .Q(StateRegOutput[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(AddRoundKeyOutput[37]), .CK(clk), .Q(StateRegOutput[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(AddRoundKeyOutput[38]), .CK(clk), .Q(StateRegOutput[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(AddRoundKeyOutput[39]), .CK(clk), .Q(StateRegOutput[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(AddRoundKeyOutput[40]), .CK(clk), .Q(StateRegOutput[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(AddRoundKeyOutput[41]), .CK(clk), .Q(StateRegOutput[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(AddRoundKeyOutput[42]), .CK(clk), .Q(StateRegOutput[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(AddRoundKeyOutput[43]), .CK(clk), .Q(StateRegOutput[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(AddRoundKeyOutput[44]), .CK(clk), .Q(StateRegOutput[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(AddRoundKeyOutput[45]), .CK(clk), .Q(StateRegOutput[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(AddRoundKeyOutput[46]), .CK(clk), .Q(StateRegOutput[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(AddRoundKeyOutput[47]), .CK(clk), .Q(StateRegOutput[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(AddRoundKeyOutput[48]), .CK(clk), .Q(StateRegOutput[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(AddRoundKeyOutput[49]), .CK(clk), .Q(StateRegOutput[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(AddRoundKeyOutput[50]), .CK(clk), .Q(StateRegOutput[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(AddRoundKeyOutput[51]), .CK(clk), .Q(StateRegOutput[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(AddRoundKeyOutput[52]), .CK(clk), .Q(StateRegOutput[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(AddRoundKeyOutput[53]), .CK(clk), .Q(StateRegOutput[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(AddRoundKeyOutput[54]), .CK(clk), .Q(StateRegOutput[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(AddRoundKeyOutput[55]), .CK(clk), .Q(StateRegOutput[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(AddRoundKeyOutput[56]), .CK(clk), .Q(StateRegOutput[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(AddRoundKeyOutput[57]), .CK(clk), .Q(StateRegOutput[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(AddRoundKeyOutput[58]), .CK(clk), .Q(StateRegOutput[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(AddRoundKeyOutput[59]), .CK(clk), .Q(StateRegOutput[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(AddRoundKeyOutput[60]), .CK(clk), .Q(StateRegOutput[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(AddRoundKeyOutput[61]), .CK(clk), .Q(StateRegOutput[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(AddRoundKeyOutput[62]), .CK(clk), .Q(StateRegOutput[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(AddRoundKeyOutput[63]), .CK(clk), .Q(StateRegOutput[63]), .QN() );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n15), .ZN(Feedback[60]) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U14 ( .A(
        StateRegOutput[1]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n10), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U13 ( .A1(
        CipherErrorVec[2]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n9), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U12 ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U9 ( .A(
        StateRegOutput[2]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n6), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U8 ( .A1(
        CipherErrorVec[1]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n5), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U7 ( .A(
        StateRegOutput[3]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n4), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U6 ( .A1(
        CipherErrorVec[0]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n3), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U5 ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n2), .B(StateRegOutput[0]), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U2 ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_U1 ( .A(CipherErrorVec[1]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_0_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n37), .ZN(Feedback[61]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U10 ( .A(
        StateRegOutput[2]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n32), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U9 ( .A1(
        CipherErrorVec[1]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U7 ( .A(
        StateRegOutput[3]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n30), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U6 ( .A1(
        CipherErrorVec[0]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U5 ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U4 ( .A(
        StateRegOutput[0]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n28), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U3 ( .A1(
        CipherErrorVec[1]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_U1 ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[2]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_1_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n15), .ZN(Feedback[62]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n8), .B(StateRegOutput[2]), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U12 ( .A1(
        CipherErrorVec[1]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n7), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U11 ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U10 ( .A(
        StateRegOutput[1]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n6), 
        .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U9 ( .A1(
        CipherErrorVec[2]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n5), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U7 ( .A(
        StateRegOutput[3]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n4), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U6 ( .A1(
        CipherErrorVec[0]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n3), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U5 ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[1]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U4 ( .A(
        StateRegOutput[0]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n2), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U2 ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_U1 ( .A(CipherErrorVec[2]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_2_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U20 ( .A(
        CipherErrorVec[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n35), .ZN(Feedback[63]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n22), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U16 ( .A1(
        StateRegOutput[3]), .A2(StateRegOutput[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U13 ( .A(
        StateRegOutput[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n36), .A2(
        StateRegOutput[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n27), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n25), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n28) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U10 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n26), .B(StateRegOutput[1]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n27) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U9 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n18), .A2(
        CipherErrorVec[2]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n26) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n21), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n25) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U7 ( .A(
        StateRegOutput[3]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n23), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n24) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U6 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n22), .A2(
        CipherErrorVec[0]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n23) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U5 ( .A1(
        CipherErrorVec[2]), .A2(CipherErrorVec[1]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n22) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U4 ( .A(
        StateRegOutput[2]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n20), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n21) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U3 ( .A1(
        CipherErrorVec[1]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n19), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n20) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U2 ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[2]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_U1 ( .A1(
        CipherErrorVec[0]), .A2(CipherErrorVec[1]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_3_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n15), .ZN(Feedback[48]) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U14 ( .A(
        StateRegOutput[5]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n10), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U13 ( .A1(
        CipherErrorVec[5]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n9), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U12 ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U9 ( .A(
        StateRegOutput[6]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n6), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U8 ( .A1(
        CipherErrorVec[4]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n5), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U7 ( .A(
        StateRegOutput[7]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n4), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U6 ( .A1(
        CipherErrorVec[3]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n3), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U5 ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n2), .B(StateRegOutput[4]), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U2 ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_U1 ( .A(CipherErrorVec[4]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_4_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n37), .ZN(Feedback[49]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U10 ( .A(
        StateRegOutput[6]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n32), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U9 ( .A1(
        CipherErrorVec[4]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U7 ( .A(
        StateRegOutput[7]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n30), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U6 ( .A1(
        CipherErrorVec[3]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U5 ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U4 ( .A(
        StateRegOutput[4]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n28), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U3 ( .A1(
        CipherErrorVec[4]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_U1 ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[5]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_5_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n15), .ZN(Feedback[50]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n8), .B(StateRegOutput[6]), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U12 ( .A1(
        CipherErrorVec[4]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n7), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U11 ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U10 ( .A(
        StateRegOutput[5]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n6), 
        .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U9 ( .A1(
        CipherErrorVec[5]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n5), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U7 ( .A(
        StateRegOutput[7]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n4), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U6 ( .A1(
        CipherErrorVec[3]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n3), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U5 ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[4]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U4 ( .A(
        StateRegOutput[4]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n2), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U2 ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_U1 ( .A(CipherErrorVec[5]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_6_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U20 ( .A(
        CipherErrorVec[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n35), .ZN(Feedback[51]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U16 ( .A1(
        StateRegOutput[7]), .A2(StateRegOutput[4]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U13 ( .A(
        StateRegOutput[7]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n36), .A2(
        StateRegOutput[4]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U9 ( .A(
        StateRegOutput[7]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n25), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n24), .A2(
        CipherErrorVec[3]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U7 ( .A1(
        CipherErrorVec[5]), .A2(CipherErrorVec[4]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U6 ( .A(
        StateRegOutput[6]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n22), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U5 ( .A1(
        CipherErrorVec[4]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U4 ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[5]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n19), .B(StateRegOutput[5]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n18), .A2(
        CipherErrorVec[5]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_U1 ( .A1(
        CipherErrorVec[3]), .A2(CipherErrorVec[4]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_7_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n15), .ZN(Feedback[52]) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U14 ( .A(
        StateRegOutput[9]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n10), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U13 ( .A1(
        CipherErrorVec[8]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n9), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U12 ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[6]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U9 ( .A(
        StateRegOutput[10]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n6), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U8 ( .A1(
        CipherErrorVec[7]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n5), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U7 ( .A(
        StateRegOutput[11]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n4), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U6 ( .A1(
        CipherErrorVec[6]), .A2(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n3), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U5 ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n2), .B(StateRegOutput[8]), 
        .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U2 ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[6]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_U1 ( .A(CipherErrorVec[7]), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_8_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n37), .ZN(Feedback[53]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U10 ( .A(
        StateRegOutput[10]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U9 ( .A1(
        CipherErrorVec[7]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U7 ( .A(
        StateRegOutput[11]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U6 ( .A1(
        CipherErrorVec[6]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U5 ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U4 ( .A(
        StateRegOutput[8]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n28), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U3 ( .A1(
        CipherErrorVec[7]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_U1 ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_9_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n15), .ZN(Feedback[54])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n8), .B(
        StateRegOutput[10]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U12 ( .A1(
        CipherErrorVec[7]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U11 ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[6]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U10 ( .A(
        StateRegOutput[9]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n6), .Z(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U9 ( .A1(
        CipherErrorVec[8]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U7 ( .A(
        StateRegOutput[11]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U6 ( .A1(
        CipherErrorVec[6]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U5 ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[7]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U4 ( .A(
        StateRegOutput[8]), .B(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n2), .ZN(SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U2 ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[6]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_U1 ( .A(
        CipherErrorVec[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_10_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U20 ( .A(
        CipherErrorVec[6]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n35), .ZN(Feedback[55])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U16 ( .A1(
        StateRegOutput[11]), .A2(StateRegOutput[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U13 ( .A(
        StateRegOutput[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n36), .A2(
        StateRegOutput[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U9 ( .A(
        StateRegOutput[11]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n24), .A2(
        CipherErrorVec[6]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U7 ( .A1(
        CipherErrorVec[8]), .A2(CipherErrorVec[7]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U6 ( .A(
        StateRegOutput[10]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U5 ( .A1(
        CipherErrorVec[7]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U4 ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n19), .B(
        StateRegOutput[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n18), .A2(
        CipherErrorVec[8]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_U1 ( .A1(
        CipherErrorVec[6]), .A2(CipherErrorVec[7]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_11_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n15), .ZN(Feedback[56])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U14 ( .A(
        StateRegOutput[13]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U13 ( .A1(
        CipherErrorVec[11]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U12 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U9 ( .A(
        StateRegOutput[14]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U8 ( .A1(
        CipherErrorVec[10]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U7 ( .A(
        StateRegOutput[15]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U6 ( .A1(
        CipherErrorVec[9]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U5 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n2), .B(
        StateRegOutput[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U2 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_U1 ( .A(
        CipherErrorVec[10]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_12_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n37), .ZN(Feedback[57])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U10 ( .A(
        StateRegOutput[14]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U9 ( .A1(
        CipherErrorVec[10]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U7 ( .A(
        StateRegOutput[15]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U6 ( .A1(
        CipherErrorVec[9]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U5 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U4 ( .A(
        StateRegOutput[12]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U3 ( .A1(
        CipherErrorVec[10]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_U1 ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_13_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n15), .ZN(Feedback[58])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n8), .B(
        StateRegOutput[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U12 ( .A1(
        CipherErrorVec[10]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U11 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U10 ( .A(
        StateRegOutput[13]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U9 ( .A1(
        CipherErrorVec[11]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U7 ( .A(
        StateRegOutput[15]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U6 ( .A1(
        CipherErrorVec[9]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U5 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[10]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U4 ( .A(
        StateRegOutput[12]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U2 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_U1 ( .A(
        CipherErrorVec[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_14_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U20 ( .A(
        CipherErrorVec[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n27), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n34), .ZN(Feedback[59])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n31), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n32), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U16 ( .A1(
        StateRegOutput[15]), .A2(StateRegOutput[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n31) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n30) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U13 ( .A(
        StateRegOutput[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n29) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n35), .A2(
        StateRegOutput[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n26), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n27) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U10 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n25), .B(
        StateRegOutput[13]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U9 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n17), .A2(
        CipherErrorVec[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n23), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U7 ( .A(
        StateRegOutput[15]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U6 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n21), .A2(
        CipherErrorVec[9]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U5 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[10]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n21) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U4 ( .A(
        StateRegOutput[14]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n19), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U3 ( .A1(
        CipherErrorVec[10]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n18), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U2 ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[11]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n18) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_U1 ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[10]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_15_n17) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n15), .ZN(Feedback[32])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U14 ( .A(
        StateRegOutput[17]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U13 ( .A1(
        CipherErrorVec[14]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U12 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U9 ( .A(
        StateRegOutput[18]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U8 ( .A1(
        CipherErrorVec[13]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U7 ( .A(
        StateRegOutput[19]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U6 ( .A1(
        CipherErrorVec[12]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U5 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n2), .B(
        StateRegOutput[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U2 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_U1 ( .A(
        CipherErrorVec[13]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_16_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n37), .ZN(Feedback[33])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U10 ( .A(
        StateRegOutput[18]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U9 ( .A1(
        CipherErrorVec[13]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U7 ( .A(
        StateRegOutput[19]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U6 ( .A1(
        CipherErrorVec[12]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U5 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U4 ( .A(
        StateRegOutput[16]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U3 ( .A1(
        CipherErrorVec[13]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_U1 ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_17_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n15), .ZN(Feedback[34])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n8), .B(
        StateRegOutput[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U12 ( .A1(
        CipherErrorVec[13]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U11 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U10 ( .A(
        StateRegOutput[17]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U9 ( .A1(
        CipherErrorVec[14]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U7 ( .A(
        StateRegOutput[19]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U6 ( .A1(
        CipherErrorVec[12]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U5 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[13]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U4 ( .A(
        StateRegOutput[16]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U2 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_U1 ( .A(
        CipherErrorVec[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_18_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U20 ( .A(
        CipherErrorVec[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n35), .ZN(Feedback[35])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U16 ( .A1(
        StateRegOutput[19]), .A2(StateRegOutput[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U13 ( .A(
        StateRegOutput[19]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n36), .A2(
        StateRegOutput[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U9 ( .A(
        StateRegOutput[19]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n24), .A2(
        CipherErrorVec[12]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U7 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[13]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U6 ( .A(
        StateRegOutput[18]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U5 ( .A1(
        CipherErrorVec[13]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U4 ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n19), .B(
        StateRegOutput[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n18), .A2(
        CipherErrorVec[14]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_U1 ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[13]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_19_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n15), .ZN(Feedback[44])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U14 ( .A(
        StateRegOutput[21]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U13 ( .A1(
        CipherErrorVec[17]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U12 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U9 ( .A(
        StateRegOutput[22]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U8 ( .A1(
        CipherErrorVec[16]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U7 ( .A(
        StateRegOutput[23]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U6 ( .A1(
        CipherErrorVec[15]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U5 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n2), .B(
        StateRegOutput[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U2 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_U1 ( .A(
        CipherErrorVec[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_20_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n37), .ZN(Feedback[45])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U10 ( .A(
        StateRegOutput[22]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U9 ( .A1(
        CipherErrorVec[16]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U7 ( .A(
        StateRegOutput[23]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U6 ( .A1(
        CipherErrorVec[15]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U5 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U4 ( .A(
        StateRegOutput[20]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U3 ( .A1(
        CipherErrorVec[16]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_U1 ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_21_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n15), .ZN(Feedback[46])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n8), .B(
        StateRegOutput[22]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U12 ( .A1(
        CipherErrorVec[16]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U11 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U10 ( .A(
        StateRegOutput[21]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U9 ( .A1(
        CipherErrorVec[17]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U7 ( .A(
        StateRegOutput[23]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U6 ( .A1(
        CipherErrorVec[15]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U5 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U4 ( .A(
        StateRegOutput[20]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U2 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_U1 ( .A(
        CipherErrorVec[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_22_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U20 ( .A(
        CipherErrorVec[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n35), .ZN(Feedback[47])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U16 ( .A1(
        StateRegOutput[23]), .A2(StateRegOutput[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U13 ( .A(
        StateRegOutput[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n36), .A2(
        StateRegOutput[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U9 ( .A(
        StateRegOutput[23]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n24), .A2(
        CipherErrorVec[15]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U7 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U6 ( .A(
        StateRegOutput[22]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U5 ( .A1(
        CipherErrorVec[16]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U4 ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n19), .B(
        StateRegOutput[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n18), .A2(
        CipherErrorVec[17]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_U1 ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[16]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_23_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n15), .ZN(Feedback[40])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U14 ( .A(
        StateRegOutput[25]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U13 ( .A1(
        CipherErrorVec[20]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U12 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U9 ( .A(
        StateRegOutput[26]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U8 ( .A1(
        CipherErrorVec[19]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U7 ( .A(
        StateRegOutput[27]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U6 ( .A1(
        CipherErrorVec[18]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U5 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n2), .B(
        StateRegOutput[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U2 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_U1 ( .A(
        CipherErrorVec[19]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_24_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n37), .ZN(Feedback[41])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U10 ( .A(
        StateRegOutput[26]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U9 ( .A1(
        CipherErrorVec[19]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U7 ( .A(
        StateRegOutput[27]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U6 ( .A1(
        CipherErrorVec[18]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U5 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U4 ( .A(
        StateRegOutput[24]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U3 ( .A1(
        CipherErrorVec[19]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_U1 ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_25_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n15), .ZN(Feedback[42])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n8), .B(
        StateRegOutput[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U12 ( .A1(
        CipherErrorVec[19]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U11 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U10 ( .A(
        StateRegOutput[25]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U9 ( .A1(
        CipherErrorVec[20]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U7 ( .A(
        StateRegOutput[27]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U6 ( .A1(
        CipherErrorVec[18]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U5 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[19]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U4 ( .A(
        StateRegOutput[24]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U2 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_U1 ( .A(
        CipherErrorVec[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_26_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U20 ( .A(
        CipherErrorVec[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n35), .ZN(Feedback[43])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U16 ( .A1(
        StateRegOutput[27]), .A2(StateRegOutput[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U13 ( .A(
        StateRegOutput[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n36), .A2(
        StateRegOutput[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U9 ( .A(
        StateRegOutput[27]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n24), .A2(
        CipherErrorVec[18]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U7 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[19]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U6 ( .A(
        StateRegOutput[26]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U5 ( .A1(
        CipherErrorVec[19]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U4 ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n19), .B(
        StateRegOutput[25]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n18), .A2(
        CipherErrorVec[20]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_U1 ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[19]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_27_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n15), .ZN(Feedback[36])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U14 ( .A(
        StateRegOutput[29]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U13 ( .A1(
        CipherErrorVec[23]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U12 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U9 ( .A(
        StateRegOutput[30]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U8 ( .A1(
        CipherErrorVec[22]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U7 ( .A(
        StateRegOutput[31]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U6 ( .A1(
        CipherErrorVec[21]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U5 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n2), .B(
        StateRegOutput[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U2 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_U1 ( .A(
        CipherErrorVec[22]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_28_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n37), .ZN(Feedback[37])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U10 ( .A(
        StateRegOutput[30]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U9 ( .A1(
        CipherErrorVec[22]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U7 ( .A(
        StateRegOutput[31]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U6 ( .A1(
        CipherErrorVec[21]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U5 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U4 ( .A(
        StateRegOutput[28]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U3 ( .A1(
        CipherErrorVec[22]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_U1 ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_29_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n15), .ZN(Feedback[38])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n8), .B(
        StateRegOutput[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U12 ( .A1(
        CipherErrorVec[22]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U11 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U10 ( .A(
        StateRegOutput[29]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U9 ( .A1(
        CipherErrorVec[23]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U7 ( .A(
        StateRegOutput[31]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U6 ( .A1(
        CipherErrorVec[21]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U5 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[22]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U4 ( .A(
        StateRegOutput[28]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U2 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_U1 ( .A(
        CipherErrorVec[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_30_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U20 ( .A(
        CipherErrorVec[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n35), .ZN(Feedback[39])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U16 ( .A1(
        StateRegOutput[31]), .A2(StateRegOutput[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U13 ( .A(
        StateRegOutput[31]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n36), .A2(
        StateRegOutput[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U9 ( .A(
        StateRegOutput[31]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n24), .A2(
        CipherErrorVec[21]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U7 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[22]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U6 ( .A(
        StateRegOutput[30]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U5 ( .A1(
        CipherErrorVec[22]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U4 ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n19), .B(
        StateRegOutput[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n18), .A2(
        CipherErrorVec[23]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_U1 ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[22]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_31_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n15), .ZN(Feedback[16])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U14 ( .A(
        StateRegOutput[33]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U13 ( .A1(
        CipherErrorVec[26]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U12 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U9 ( .A(
        StateRegOutput[34]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U8 ( .A1(
        CipherErrorVec[25]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U7 ( .A(
        StateRegOutput[35]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U6 ( .A1(
        CipherErrorVec[24]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U5 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n2), .B(
        StateRegOutput[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U2 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_U1 ( .A(
        CipherErrorVec[25]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_32_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n37), .ZN(Feedback[17])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U10 ( .A(
        StateRegOutput[34]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U9 ( .A1(
        CipherErrorVec[25]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U7 ( .A(
        StateRegOutput[35]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U6 ( .A1(
        CipherErrorVec[24]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U5 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U4 ( .A(
        StateRegOutput[32]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U3 ( .A1(
        CipherErrorVec[25]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_U1 ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_33_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n15), .ZN(Feedback[18])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n8), .B(
        StateRegOutput[34]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U12 ( .A1(
        CipherErrorVec[25]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U11 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U10 ( .A(
        StateRegOutput[33]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U9 ( .A1(
        CipherErrorVec[26]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U7 ( .A(
        StateRegOutput[35]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U6 ( .A1(
        CipherErrorVec[24]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U5 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[25]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U4 ( .A(
        StateRegOutput[32]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U2 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_U1 ( .A(
        CipherErrorVec[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_34_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U20 ( .A(
        CipherErrorVec[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n35), .ZN(Feedback[19])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U16 ( .A1(
        StateRegOutput[35]), .A2(StateRegOutput[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U13 ( .A(
        StateRegOutput[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n36), .A2(
        StateRegOutput[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U9 ( .A(
        StateRegOutput[35]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n24), .A2(
        CipherErrorVec[24]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U7 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[25]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U6 ( .A(
        StateRegOutput[34]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U5 ( .A1(
        CipherErrorVec[25]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U4 ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n19), .B(
        StateRegOutput[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n18), .A2(
        CipherErrorVec[26]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_U1 ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[25]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_35_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n15), .ZN(Feedback[28])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U14 ( .A(
        StateRegOutput[37]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U13 ( .A1(
        CipherErrorVec[29]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U12 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U9 ( .A(
        StateRegOutput[38]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U8 ( .A1(
        CipherErrorVec[28]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U7 ( .A(
        StateRegOutput[39]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U6 ( .A1(
        CipherErrorVec[27]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U5 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n2), .B(
        StateRegOutput[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U2 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_U1 ( .A(
        CipherErrorVec[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_36_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n37), .ZN(Feedback[29])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U10 ( .A(
        StateRegOutput[38]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U9 ( .A1(
        CipherErrorVec[28]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U7 ( .A(
        StateRegOutput[39]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U6 ( .A1(
        CipherErrorVec[27]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U5 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U4 ( .A(
        StateRegOutput[36]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U3 ( .A1(
        CipherErrorVec[28]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_U1 ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_37_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n15), .ZN(Feedback[30])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n8), .B(
        StateRegOutput[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U12 ( .A1(
        CipherErrorVec[28]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U11 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U10 ( .A(
        StateRegOutput[37]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U9 ( .A1(
        CipherErrorVec[29]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U7 ( .A(
        StateRegOutput[39]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U6 ( .A1(
        CipherErrorVec[27]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U5 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U4 ( .A(
        StateRegOutput[36]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U2 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_U1 ( .A(
        CipherErrorVec[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_38_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U20 ( .A(
        CipherErrorVec[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n35), .ZN(Feedback[31])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U16 ( .A1(
        StateRegOutput[39]), .A2(StateRegOutput[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U13 ( .A(
        StateRegOutput[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n36), .A2(
        StateRegOutput[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U9 ( .A(
        StateRegOutput[39]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n24), .A2(
        CipherErrorVec[27]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U7 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U6 ( .A(
        StateRegOutput[38]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U5 ( .A1(
        CipherErrorVec[28]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U4 ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n19), .B(
        StateRegOutput[37]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n18), .A2(
        CipherErrorVec[29]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_U1 ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[28]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_39_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n15), .ZN(Feedback[24])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U14 ( .A(
        StateRegOutput[41]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U13 ( .A1(
        CipherErrorVec[32]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U12 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U9 ( .A(
        StateRegOutput[42]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U8 ( .A1(
        CipherErrorVec[31]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U7 ( .A(
        StateRegOutput[43]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U6 ( .A1(
        CipherErrorVec[30]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U5 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n2), .B(
        StateRegOutput[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U2 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_U1 ( .A(
        CipherErrorVec[31]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_40_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n37), .ZN(Feedback[25])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U10 ( .A(
        StateRegOutput[42]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U9 ( .A1(
        CipherErrorVec[31]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U7 ( .A(
        StateRegOutput[43]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U6 ( .A1(
        CipherErrorVec[30]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U5 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U4 ( .A(
        StateRegOutput[40]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U3 ( .A1(
        CipherErrorVec[31]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_U1 ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_41_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n15), .ZN(Feedback[26])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n8), .B(
        StateRegOutput[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U12 ( .A1(
        CipherErrorVec[31]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U11 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U10 ( .A(
        StateRegOutput[41]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U9 ( .A1(
        CipherErrorVec[32]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U7 ( .A(
        StateRegOutput[43]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U6 ( .A1(
        CipherErrorVec[30]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U5 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[31]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U4 ( .A(
        StateRegOutput[40]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U2 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_U1 ( .A(
        CipherErrorVec[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_42_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U20 ( .A(
        CipherErrorVec[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n35), .ZN(Feedback[27])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U16 ( .A1(
        StateRegOutput[43]), .A2(StateRegOutput[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U13 ( .A(
        StateRegOutput[43]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n36), .A2(
        StateRegOutput[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U9 ( .A(
        StateRegOutput[43]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n24), .A2(
        CipherErrorVec[30]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U7 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[31]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U6 ( .A(
        StateRegOutput[42]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U5 ( .A1(
        CipherErrorVec[31]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U4 ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n19), .B(
        StateRegOutput[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n18), .A2(
        CipherErrorVec[32]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_U1 ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[31]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_43_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n15), .ZN(Feedback[20])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U14 ( .A(
        StateRegOutput[45]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U13 ( .A1(
        CipherErrorVec[35]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U12 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U9 ( .A(
        StateRegOutput[46]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U8 ( .A1(
        CipherErrorVec[34]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U7 ( .A(
        StateRegOutput[47]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U6 ( .A1(
        CipherErrorVec[33]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U5 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n2), .B(
        StateRegOutput[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U2 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_U1 ( .A(
        CipherErrorVec[34]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_44_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n37), .ZN(Feedback[21])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U10 ( .A(
        StateRegOutput[46]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U9 ( .A1(
        CipherErrorVec[34]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U7 ( .A(
        StateRegOutput[47]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U6 ( .A1(
        CipherErrorVec[33]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U5 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U4 ( .A(
        StateRegOutput[44]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U3 ( .A1(
        CipherErrorVec[34]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_U1 ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_45_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n15), .ZN(Feedback[22])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n8), .B(
        StateRegOutput[46]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U12 ( .A1(
        CipherErrorVec[34]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U11 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U10 ( .A(
        StateRegOutput[45]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U9 ( .A1(
        CipherErrorVec[35]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U7 ( .A(
        StateRegOutput[47]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U6 ( .A1(
        CipherErrorVec[33]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U5 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[34]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U4 ( .A(
        StateRegOutput[44]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U2 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_U1 ( .A(
        CipherErrorVec[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_46_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U20 ( .A(
        CipherErrorVec[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n35), .ZN(Feedback[23])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U16 ( .A1(
        StateRegOutput[47]), .A2(StateRegOutput[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U13 ( .A(
        StateRegOutput[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n36), .A2(
        StateRegOutput[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U9 ( .A(
        StateRegOutput[47]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n24), .A2(
        CipherErrorVec[33]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U7 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[34]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U6 ( .A(
        StateRegOutput[46]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U5 ( .A1(
        CipherErrorVec[34]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U4 ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n19), .B(
        StateRegOutput[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n18), .A2(
        CipherErrorVec[35]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_U1 ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[34]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_47_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n15), .ZN(Feedback[4]) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U14 ( .A(
        StateRegOutput[49]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U13 ( .A1(
        CipherErrorVec[38]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U12 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U9 ( .A(
        StateRegOutput[50]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U8 ( .A1(
        CipherErrorVec[37]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U7 ( .A(
        StateRegOutput[51]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U6 ( .A1(
        CipherErrorVec[36]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U5 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n2), .B(
        StateRegOutput[48]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U2 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_U1 ( .A(
        CipherErrorVec[37]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_48_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n37), .ZN(Feedback[5]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U10 ( .A(
        StateRegOutput[50]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U9 ( .A1(
        CipherErrorVec[37]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U7 ( .A(
        StateRegOutput[51]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U6 ( .A1(
        CipherErrorVec[36]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U5 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U4 ( .A(
        StateRegOutput[48]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U3 ( .A1(
        CipherErrorVec[37]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_U1 ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_49_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n15), .ZN(Feedback[6]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n8), .B(
        StateRegOutput[50]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U12 ( .A1(
        CipherErrorVec[37]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U11 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U10 ( .A(
        StateRegOutput[49]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U9 ( .A1(
        CipherErrorVec[38]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U7 ( .A(
        StateRegOutput[51]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U6 ( .A1(
        CipherErrorVec[36]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U5 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[37]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U4 ( .A(
        StateRegOutput[48]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U2 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_U1 ( .A(
        CipherErrorVec[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_50_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U20 ( .A(
        CipherErrorVec[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n35), .ZN(Feedback[7]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U16 ( .A1(
        StateRegOutput[51]), .A2(StateRegOutput[48]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U13 ( .A(
        StateRegOutput[51]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n36), .A2(
        StateRegOutput[48]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U9 ( .A(
        StateRegOutput[51]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n24), .A2(
        CipherErrorVec[36]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U7 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[37]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U6 ( .A(
        StateRegOutput[50]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U5 ( .A1(
        CipherErrorVec[37]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U4 ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n19), .B(
        StateRegOutput[49]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n18), .A2(
        CipherErrorVec[38]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_U1 ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[37]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_51_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n15), .ZN(Feedback[8]) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U14 ( .A(
        StateRegOutput[53]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U13 ( .A1(
        CipherErrorVec[41]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U12 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U9 ( .A(
        StateRegOutput[54]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U8 ( .A1(
        CipherErrorVec[40]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U7 ( .A(
        StateRegOutput[55]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U6 ( .A1(
        CipherErrorVec[39]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U5 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n2), .B(
        StateRegOutput[52]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U2 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_U1 ( .A(
        CipherErrorVec[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_52_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n37), .ZN(Feedback[9]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U10 ( .A(
        StateRegOutput[54]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U9 ( .A1(
        CipherErrorVec[40]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U7 ( .A(
        StateRegOutput[55]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U6 ( .A1(
        CipherErrorVec[39]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U5 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U4 ( .A(
        StateRegOutput[52]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U3 ( .A1(
        CipherErrorVec[40]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_U1 ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_53_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n15), .ZN(Feedback[10])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n8), .B(
        StateRegOutput[54]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U12 ( .A1(
        CipherErrorVec[40]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U11 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U10 ( .A(
        StateRegOutput[53]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U9 ( .A1(
        CipherErrorVec[41]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U7 ( .A(
        StateRegOutput[55]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U6 ( .A1(
        CipherErrorVec[39]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U5 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U4 ( .A(
        StateRegOutput[52]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U2 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_U1 ( .A(
        CipherErrorVec[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_54_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U20 ( .A(
        CipherErrorVec[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n35), .ZN(Feedback[11])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U16 ( .A1(
        StateRegOutput[55]), .A2(StateRegOutput[52]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U13 ( .A(
        StateRegOutput[55]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n36), .A2(
        StateRegOutput[52]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U9 ( .A(
        StateRegOutput[55]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n24), .A2(
        CipherErrorVec[39]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U7 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U6 ( .A(
        StateRegOutput[54]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U5 ( .A1(
        CipherErrorVec[40]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U4 ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n19), .B(
        StateRegOutput[53]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n18), .A2(
        CipherErrorVec[41]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_U1 ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[40]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_55_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n15), .ZN(Feedback[12])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U14 ( .A(
        StateRegOutput[57]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U13 ( .A1(
        CipherErrorVec[44]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U12 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U9 ( .A(
        StateRegOutput[58]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U8 ( .A1(
        CipherErrorVec[43]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U7 ( .A(
        StateRegOutput[59]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U6 ( .A1(
        CipherErrorVec[42]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U5 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n2), .B(
        StateRegOutput[56]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U2 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_U1 ( .A(
        CipherErrorVec[43]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_56_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n37), .ZN(Feedback[13])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U10 ( .A(
        StateRegOutput[58]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U9 ( .A1(
        CipherErrorVec[43]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U7 ( .A(
        StateRegOutput[59]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U6 ( .A1(
        CipherErrorVec[42]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U5 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U4 ( .A(
        StateRegOutput[56]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U3 ( .A1(
        CipherErrorVec[43]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_U1 ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_57_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n15), .ZN(Feedback[14])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n8), .B(
        StateRegOutput[58]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U12 ( .A1(
        CipherErrorVec[43]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U11 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U10 ( .A(
        StateRegOutput[57]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U9 ( .A1(
        CipherErrorVec[44]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U7 ( .A(
        StateRegOutput[59]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U6 ( .A1(
        CipherErrorVec[42]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U5 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[43]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U4 ( .A(
        StateRegOutput[56]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U2 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_U1 ( .A(
        CipherErrorVec[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_58_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U20 ( .A(
        CipherErrorVec[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n35), .ZN(Feedback[15])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U16 ( .A1(
        StateRegOutput[59]), .A2(StateRegOutput[56]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U13 ( .A(
        StateRegOutput[59]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n36), .A2(
        StateRegOutput[56]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U9 ( .A(
        StateRegOutput[59]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n24), .A2(
        CipherErrorVec[42]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U7 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[43]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U6 ( .A(
        StateRegOutput[58]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U5 ( .A1(
        CipherErrorVec[43]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U4 ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n19), .B(
        StateRegOutput[57]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n18), .A2(
        CipherErrorVec[44]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_U1 ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[43]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_59_n18) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n15), .ZN(Feedback[0]) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n15) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n16) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U14 ( .A(
        StateRegOutput[61]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n10), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n11) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U13 ( .A1(
        CipherErrorVec[47]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n10) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U12 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n8), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n12) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n13), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n14), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n7) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U9 ( .A(
        StateRegOutput[62]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n6), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U8 ( .A1(
        CipherErrorVec[46]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n6) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U7 ( .A(
        StateRegOutput[63]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n13) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U6 ( .A1(
        CipherErrorVec[45]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U5 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U4 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n2), .B(
        StateRegOutput[60]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n8) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U2 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_U1 ( .A(
        CipherErrorVec[46]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_60_n1) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U13 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n38), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n37), .ZN(Feedback[1]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n37) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n34), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n33), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n38) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U10 ( .A(
        StateRegOutput[62]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n32), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U9 ( .A1(
        CipherErrorVec[46]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n32) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n35), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n34) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U7 ( .A(
        StateRegOutput[63]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n35) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U6 ( .A1(
        CipherErrorVec[45]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n29), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n30) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U5 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n29) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U4 ( .A(
        StateRegOutput[60]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n28), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U3 ( .A1(
        CipherErrorVec[46]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n28) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U2 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n27) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_U1 ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_61_n31) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U17 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n16), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n15), .ZN(Feedback[2]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U16 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n14), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n13), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n15) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n12), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n11), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n13) );
  OR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n11) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U13 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n8), .B(
        StateRegOutput[62]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n12) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U12 ( .A1(
        CipherErrorVec[46]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n7), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n8) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U11 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n7) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U10 ( .A(
        StateRegOutput[61]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n6), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n14) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U9 ( .A1(
        CipherErrorVec[47]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n6) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n10), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n9), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n16) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U7 ( .A(
        StateRegOutput[63]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n4), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n9) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U6 ( .A1(
        CipherErrorVec[45]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n3), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n4) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U5 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[46]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n3) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U4 ( .A(
        StateRegOutput[60]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n2), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n10) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U3 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n1), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n5), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n2) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U2 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n5) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_U1 ( .A(
        CipherErrorVec[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_62_n1) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U20 ( .A(
        CipherErrorVec[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U19 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n28), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n35), .ZN(Feedback[3]) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U18 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n32), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n34), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n35) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U17 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n33), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n24), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n34) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U16 ( .A1(
        StateRegOutput[63]), .A2(StateRegOutput[60]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n33) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U15 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n29), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n31), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n32) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U14 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n30), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n31) );
  INV_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U13 ( .A(
        StateRegOutput[63]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n30) );
  AND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U12 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n36), .A2(
        StateRegOutput[60]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n29) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U11 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n20), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n27), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n28) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U10 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n23), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n26), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n27) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U9 ( .A(
        StateRegOutput[63]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n25), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n26) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U8 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n24), .A2(
        CipherErrorVec[45]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n25) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U7 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[46]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n24) );
  XOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U6 ( .A(
        StateRegOutput[62]), .B(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n22), .Z(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n23) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U5 ( .A1(
        CipherErrorVec[46]), .A2(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n21), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n22) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U4 ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n21) );
  XNOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U3 ( .A(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n19), .B(
        StateRegOutput[61]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n20) );
  NOR2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U2 ( .A1(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n18), .A2(
        CipherErrorVec[47]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n19) );
  NAND2_X1 SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_U1 ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[46]), .ZN(
        SD1_Xor_Sbox_Inst_SD1_Xor_FMulti_bit_inst_63_n18) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n3), .B(Input[2]), .ZN(
        Red_MCOutput[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Input[0]), .B(Input[1]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_1_n3), .B(Input[3]), .ZN(
        Red_MCOutput[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U1 ( .A(Input[0]), .B(Input[1]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_2_n3), .B(Input[3]), .ZN(
        Red_MCOutput[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U1 ( .A(Input[0]), .B(Input[2]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n3), .B(Input[6]), .ZN(
        Red_MCOutput[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Input[4]), .B(Input[5]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_1_n3), .B(Input[7]), .ZN(
        Red_MCOutput[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U1 ( .A(Input[4]), .B(Input[5]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_2_n3), .B(Input[7]), .ZN(
        Red_MCOutput[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U1 ( .A(Input[4]), .B(Input[6]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n3), .B(Input[10]), .ZN(
        Red_MCOutput[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Input[8]), .B(Input[9]), 
        .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_1_n3), .B(Input[11]), .ZN(
        Red_MCOutput[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U1 ( .A(Input[8]), .B(Input[9]), 
        .ZN(Red_PlaintextInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_2_n3), .B(Input[11]), .ZN(
        Red_MCOutput[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U1 ( .A(Input[8]), .B(Input[10]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n3), .B(Input[14]), .ZN(
        Red_MCOutput[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Input[12]), .B(
        Input[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_1_n3), .B(Input[15]), .ZN(
        Red_MCOutput[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U1 ( .A(Input[12]), .B(
        Input[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_2_n3), .B(Input[15]), .ZN(
        Red_MCOutput[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U1 ( .A(Input[12]), .B(
        Input[14]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n3), .B(Input[18]), .ZN(
        Red_MCOutput[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Input[16]), .B(
        Input[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_1_n3), .B(Input[19]), .ZN(
        Red_MCOutput[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U1 ( .A(Input[16]), .B(
        Input[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_2_n3), .B(Input[19]), .ZN(
        Red_MCOutput[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U1 ( .A(Input[16]), .B(
        Input[18]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n3), .B(Input[22]), .ZN(
        Red_MCOutput[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Input[20]), .B(
        Input[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_1_n3), .B(Input[23]), .ZN(
        Red_MCOutput[16]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U1 ( .A(Input[20]), .B(
        Input[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_2_n3), .B(Input[23]), .ZN(
        Red_MCOutput[17]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U1 ( .A(Input[20]), .B(
        Input[22]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n3), .B(Input[26]), .ZN(
        Red_MCOutput[18]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Input[24]), .B(
        Input[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_1_n3), .B(Input[27]), .ZN(
        Red_MCOutput[19]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U1 ( .A(Input[24]), .B(
        Input[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_2_n3), .B(Input[27]), .ZN(
        Red_MCOutput[20]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U1 ( .A(Input[24]), .B(
        Input[26]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n3), .B(Input[30]), .ZN(
        Red_MCOutput[21]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Input[28]), .B(
        Input[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_1_n3), .B(Input[31]), .ZN(
        Red_MCOutput[22]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U1 ( .A(Input[28]), .B(
        Input[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_2_n3), .B(Input[31]), .ZN(
        Red_MCOutput[23]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U1 ( .A(Input[28]), .B(
        Input[30]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n3), .B(Input[34]), .ZN(
        Red_Input[24]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Input[32]), .B(
        Input[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_1_n3), .B(Input[35]), .ZN(
        Red_Input[25]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U1 ( .A(Input[32]), .B(
        Input[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_2_n3), .B(Input[35]), .ZN(
        Red_Input[26]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U1 ( .A(Input[32]), .B(
        Input[34]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n3), .B(Input[38]), .ZN(
        Red_Input[27]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Input[36]), .B(
        Input[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_1_n3), .B(Input[39]), .ZN(
        Red_Input[28]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U1 ( .A(Input[36]), .B(
        Input[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_2_n3), .B(Input[39]), .ZN(
        Red_Input[29]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U1 ( .A(Input[36]), .B(
        Input[38]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n3), .B(Input[42]), .ZN(
        Red_Input[30]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Input[40]), .B(
        Input[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_1_n3), .B(Input[43]), .ZN(
        Red_Input[31]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U1 ( .A(Input[40]), .B(
        Input[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_2_n3), .B(Input[43]), .ZN(
        Red_Input[32]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U1 ( .A(Input[40]), .B(
        Input[42]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n3), .B(Input[46]), .ZN(
        Red_Input[33]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Input[44]), .B(
        Input[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_1_n3), .B(Input[47]), .ZN(
        Red_Input[34]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U1 ( .A(Input[44]), .B(
        Input[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_2_n3), .B(Input[47]), .ZN(
        Red_Input[35]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U1 ( .A(Input[44]), .B(
        Input[46]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n3), .B(Input[50]), .ZN(
        Red_Input[36]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Input[48]), .B(
        Input[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_1_n3), .B(Input[51]), .ZN(
        Red_Input[37]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U1 ( .A(Input[48]), .B(
        Input[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_2_n3), .B(Input[51]), .ZN(
        Red_Input[38]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U1 ( .A(Input[48]), .B(
        Input[50]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n3), .B(Input[54]), .ZN(
        Red_Input[39]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Input[52]), .B(
        Input[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_1_n3), .B(Input[55]), .ZN(
        Red_Input[40]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U1 ( .A(Input[52]), .B(
        Input[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_2_n3), .B(Input[55]), .ZN(
        Red_Input[41]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U1 ( .A(Input[52]), .B(
        Input[54]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n3), .B(Input[58]), .ZN(
        Red_Input[42]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Input[56]), .B(
        Input[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_1_n3), .B(Input[59]), .ZN(
        Red_Input[43]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U1 ( .A(Input[56]), .B(
        Input[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_2_n3), .B(Input[59]), .ZN(
        Red_Input[44]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U1 ( .A(Input[56]), .B(
        Input[58]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n3), .B(Input[62]), .ZN(
        Red_Input[45]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Input[60]), .B(
        Input[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_1_n3), .B(Input[63]), .ZN(
        Red_Input[46]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U1 ( .A(Input[60]), .B(
        Input[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_2_n3), .B(Input[63]), .ZN(
        Red_Input[47]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U1 ( .A(Input[60]), .B(
        Input[62]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_2_n3) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U2 ( .A(Red_MCInst_XOR_r0_Inst_0_n5), .B(
        Red_MCOutput[12]), .ZN(Red_MCOutput[36]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U1 ( .A(Red_MCOutput[0]), .B(Red_Input[36]), .ZN(Red_MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_0_U1 ( .A(Red_Input[24]), .B(Red_MCOutput[0]), 
        .Z(Red_MCOutput[24]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U2 ( .A(Red_MCInst_XOR_r0_Inst_1_n5), .B(
        Red_MCOutput[13]), .ZN(Red_MCOutput[37]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U1 ( .A(Red_MCOutput[1]), .B(Red_Input[37]), .ZN(Red_MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_1_U1 ( .A(Red_Input[25]), .B(Red_MCOutput[1]), 
        .Z(Red_MCOutput[25]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U2 ( .A(Red_MCInst_XOR_r0_Inst_2_n5), .B(
        Red_MCOutput[14]), .ZN(Red_MCOutput[38]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U1 ( .A(Red_MCOutput[2]), .B(Red_Input[38]), .ZN(Red_MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_2_U1 ( .A(Red_Input[26]), .B(Red_MCOutput[2]), 
        .Z(Red_MCOutput[26]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U2 ( .A(Red_MCInst_XOR_r0_Inst_3_n5), .B(
        Red_MCOutput[15]), .ZN(Red_MCOutput[39]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U1 ( .A(Red_MCOutput[3]), .B(Red_Input[39]), .ZN(Red_MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_3_U1 ( .A(Red_Input[27]), .B(Red_MCOutput[3]), 
        .Z(Red_MCOutput[27]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_4_U2 ( .A(Red_MCInst_XOR_r0_Inst_4_n5), .B(
        Red_MCOutput[16]), .ZN(Red_MCOutput[40]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_4_U1 ( .A(Red_MCOutput[4]), .B(Red_Input[40]), .ZN(Red_MCInst_XOR_r0_Inst_4_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_4_U1 ( .A(Red_Input[28]), .B(Red_MCOutput[4]), 
        .Z(Red_MCOutput[28]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_5_U2 ( .A(Red_MCInst_XOR_r0_Inst_5_n5), .B(
        Red_MCOutput[17]), .ZN(Red_MCOutput[41]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_5_U1 ( .A(Red_MCOutput[5]), .B(Red_Input[41]), .ZN(Red_MCInst_XOR_r0_Inst_5_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_5_U1 ( .A(Red_Input[29]), .B(Red_MCOutput[5]), 
        .Z(Red_MCOutput[29]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_6_U2 ( .A(Red_MCInst_XOR_r0_Inst_6_n5), .B(
        Red_MCOutput[18]), .ZN(Red_MCOutput[42]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_6_U1 ( .A(Red_MCOutput[6]), .B(Red_Input[42]), .ZN(Red_MCInst_XOR_r0_Inst_6_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_6_U1 ( .A(Red_Input[30]), .B(Red_MCOutput[6]), 
        .Z(Red_MCOutput[30]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_7_U2 ( .A(Red_MCInst_XOR_r0_Inst_7_n5), .B(
        Red_MCOutput[19]), .ZN(Red_MCOutput[43]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_7_U1 ( .A(Red_MCOutput[7]), .B(Red_Input[43]), .ZN(Red_MCInst_XOR_r0_Inst_7_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_7_U1 ( .A(Red_Input[31]), .B(Red_MCOutput[7]), 
        .Z(Red_MCOutput[31]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_8_U2 ( .A(Red_MCInst_XOR_r0_Inst_8_n5), .B(
        Red_MCOutput[20]), .ZN(Red_MCOutput[44]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_8_U1 ( .A(Red_MCOutput[8]), .B(Red_Input[44]), .ZN(Red_MCInst_XOR_r0_Inst_8_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_8_U1 ( .A(Red_Input[32]), .B(Red_MCOutput[8]), 
        .Z(Red_MCOutput[32]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_9_U2 ( .A(Red_MCInst_XOR_r0_Inst_9_n5), .B(
        Red_MCOutput[21]), .ZN(Red_MCOutput[45]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_9_U1 ( .A(Red_MCOutput[9]), .B(Red_Input[45]), .ZN(Red_MCInst_XOR_r0_Inst_9_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_9_U1 ( .A(Red_Input[33]), .B(Red_MCOutput[9]), 
        .Z(Red_MCOutput[33]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_10_U2 ( .A(Red_MCInst_XOR_r0_Inst_10_n5), 
        .B(Red_MCOutput[22]), .ZN(Red_MCOutput[46]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_10_U1 ( .A(Red_MCOutput[10]), .B(
        Red_Input[46]), .ZN(Red_MCInst_XOR_r0_Inst_10_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_10_U1 ( .A(Red_Input[34]), .B(
        Red_MCOutput[10]), .Z(Red_MCOutput[34]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_11_U2 ( .A(Red_MCInst_XOR_r0_Inst_11_n5), 
        .B(Red_MCOutput[23]), .ZN(Red_MCOutput[47]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_11_U1 ( .A(Red_MCOutput[11]), .B(
        Red_Input[47]), .ZN(Red_MCInst_XOR_r0_Inst_11_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_11_U1 ( .A(Red_Input[35]), .B(
        Red_MCOutput[11]), .Z(Red_MCOutput[35]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_0_U1 ( .A(Red_MCOutput[36]), .B(Red_K1[36]), 
        .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_1_U1 ( .A(Red_MCOutput[37]), .B(Red_K1[37]), 
        .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_2_U1 ( .A(Red_MCOutput[38]), .B(Red_K1[38]), 
        .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_0_U1 ( .A(Red_MCOutput[39]), .B(Red_K1[39]), 
        .Z(Red_AddRoundKeyOutput[39]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_1_U1 ( .A(Red_MCOutput[40]), .B(Red_K1[40]), 
        .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_2_U1 ( .A(Red_MCOutput[41]), .B(Red_K1[41]), 
        .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_0_U1 ( .A(Red_MCOutput[42]), .B(Red_K1[42]), 
        .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_1_U1 ( .A(Red_MCOutput[43]), .B(Red_K1[43]), 
        .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_2_U1 ( .A(Red_MCOutput[44]), .B(Red_K1[44]), 
        .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_0_U1 ( .A(Red_MCOutput[45]), .B(Red_K1[45]), 
        .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_1_U1 ( .A(Red_MCOutput[46]), .B(Red_K1[46]), 
        .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_2_U1 ( .A(Red_MCOutput[47]), .B(Red_K1[47]), 
        .Z(Red_AddRoundKeyOutput[47]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U1 ( .A(Red_MCOutput[30]), .B(
        Red_K1[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_1_U1 ( .A(Red_MCOutput[31]), .B(
        Red_K1[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_2_U1 ( .A(Red_MCOutput[32]), .B(
        Red_K1[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U1 ( .A(Red_MCOutput[33]), .B(
        Red_K1[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_1_U1 ( .A(Red_MCOutput[34]), .B(
        Red_K1[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_2_U1 ( .A(Red_MCOutput[35]), .B(
        Red_K1[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_0_U1 ( .A(Red_MCOutput[0]), .B(Red_K1[0]), 
        .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_1_U1 ( .A(Red_MCOutput[1]), .B(Red_K1[1]), 
        .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_2_U1 ( .A(Red_MCOutput[2]), .B(Red_K1[2]), 
        .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_0_U1 ( .A(Red_MCOutput[3]), .B(Red_K1[3]), 
        .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_1_U1 ( .A(Red_MCOutput[4]), .B(Red_K1[4]), 
        .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_2_U1 ( .A(Red_MCOutput[5]), .B(Red_K1[5]), 
        .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_0_U1 ( .A(Red_MCOutput[6]), .B(Red_K1[6]), 
        .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_1_U1 ( .A(Red_MCOutput[7]), .B(Red_K1[7]), 
        .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_2_U1 ( .A(Red_MCOutput[8]), .B(Red_K1[8]), 
        .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_0_U1 ( .A(Red_MCOutput[9]), .B(Red_K1[9]), 
        .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_1_U1 ( .A(Red_MCOutput[10]), .B(Red_K1[10]), 
        .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_2_U1 ( .A(Red_MCOutput[11]), .B(Red_K1[11]), 
        .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_0_U1 ( .A(Red_MCOutput[12]), .B(Red_K1[12]), 
        .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_1_U1 ( .A(Red_MCOutput[13]), .B(Red_K1[13]), 
        .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_2_U1 ( .A(Red_MCOutput[14]), .B(Red_K1[14]), 
        .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_0_U1 ( .A(Red_MCOutput[15]), .B(Red_K1[15]), 
        .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_1_U1 ( .A(Red_MCOutput[16]), .B(Red_K1[16]), 
        .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_2_U1 ( .A(Red_MCOutput[17]), .B(Red_K1[17]), 
        .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_0_U1 ( .A(Red_MCOutput[18]), .B(Red_K1[18]), 
        .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_1_U1 ( .A(Red_MCOutput[19]), .B(Red_K1[19]), 
        .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_2_U1 ( .A(Red_MCOutput[20]), .B(Red_K1[20]), 
        .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_0_U1 ( .A(Red_MCOutput[21]), .B(Red_K1[21]), 
        .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_1_U1 ( .A(Red_MCOutput[22]), .B(Red_K1[22]), 
        .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_2_U1 ( .A(Red_MCOutput[23]), .B(Red_K1[23]), 
        .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_0_U1 ( .A(Red_MCOutput[24]), .B(Red_K1[24]), 
        .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_1_U1 ( .A(Red_MCOutput[25]), .B(Red_K1[25]), 
        .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_2_U1 ( .A(Red_MCOutput[26]), .B(Red_K1[26]), 
        .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_0_U1 ( .A(Red_MCOutput[27]), .B(Red_K1[27]), 
        .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_1_U1 ( .A(Red_MCOutput[28]), .B(Red_K1[28]), 
        .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_2_U1 ( .A(Red_MCOutput[29]), .B(Red_K1[29]), 
        .Z(Red_AddRoundKeyOutput[29]) );
  DFF_X1 Red_StateReg_s_current_state_reg_0_ ( .D(Red_AddRoundKeyOutput[0]), 
        .CK(clk), .Q(Red_StateRegOutput[0]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_1_ ( .D(Red_AddRoundKeyOutput[1]), 
        .CK(clk), .Q(Red_StateRegOutput[1]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_2_ ( .D(Red_AddRoundKeyOutput[2]), 
        .CK(clk), .Q(Red_StateRegOutput[2]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_3_ ( .D(Red_AddRoundKeyOutput[3]), 
        .CK(clk), .Q(Red_StateRegOutput[3]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_4_ ( .D(Red_AddRoundKeyOutput[4]), 
        .CK(clk), .Q(Red_StateRegOutput[4]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_5_ ( .D(Red_AddRoundKeyOutput[5]), 
        .CK(clk), .Q(Red_StateRegOutput[5]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_6_ ( .D(Red_AddRoundKeyOutput[6]), 
        .CK(clk), .Q(Red_StateRegOutput[6]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_7_ ( .D(Red_AddRoundKeyOutput[7]), 
        .CK(clk), .Q(Red_StateRegOutput[7]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_8_ ( .D(Red_AddRoundKeyOutput[8]), 
        .CK(clk), .Q(Red_StateRegOutput[8]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_9_ ( .D(Red_AddRoundKeyOutput[9]), 
        .CK(clk), .Q(Red_StateRegOutput[9]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_10_ ( .D(Red_AddRoundKeyOutput[10]), 
        .CK(clk), .Q(Red_StateRegOutput[10]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_11_ ( .D(Red_AddRoundKeyOutput[11]), 
        .CK(clk), .Q(Red_StateRegOutput[11]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_12_ ( .D(Red_AddRoundKeyOutput[12]), 
        .CK(clk), .Q(Red_StateRegOutput[12]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_13_ ( .D(Red_AddRoundKeyOutput[13]), 
        .CK(clk), .Q(Red_StateRegOutput[13]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_14_ ( .D(Red_AddRoundKeyOutput[14]), 
        .CK(clk), .Q(Red_StateRegOutput[14]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_15_ ( .D(Red_AddRoundKeyOutput[15]), 
        .CK(clk), .Q(Red_StateRegOutput[15]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_16_ ( .D(Red_AddRoundKeyOutput[16]), 
        .CK(clk), .Q(Red_StateRegOutput[16]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_17_ ( .D(Red_AddRoundKeyOutput[17]), 
        .CK(clk), .Q(Red_StateRegOutput[17]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_18_ ( .D(Red_AddRoundKeyOutput[18]), 
        .CK(clk), .Q(Red_StateRegOutput[18]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_19_ ( .D(Red_AddRoundKeyOutput[19]), 
        .CK(clk), .Q(Red_StateRegOutput[19]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_20_ ( .D(Red_AddRoundKeyOutput[20]), 
        .CK(clk), .Q(Red_StateRegOutput[20]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_21_ ( .D(Red_AddRoundKeyOutput[21]), 
        .CK(clk), .Q(Red_StateRegOutput[21]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_22_ ( .D(Red_AddRoundKeyOutput[22]), 
        .CK(clk), .Q(Red_StateRegOutput[22]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_23_ ( .D(Red_AddRoundKeyOutput[23]), 
        .CK(clk), .Q(Red_StateRegOutput[23]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_24_ ( .D(Red_AddRoundKeyOutput[24]), 
        .CK(clk), .Q(Red_StateRegOutput[24]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_25_ ( .D(Red_AddRoundKeyOutput[25]), 
        .CK(clk), .Q(Red_StateRegOutput[25]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_26_ ( .D(Red_AddRoundKeyOutput[26]), 
        .CK(clk), .Q(Red_StateRegOutput[26]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_27_ ( .D(Red_AddRoundKeyOutput[27]), 
        .CK(clk), .Q(Red_StateRegOutput[27]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_28_ ( .D(Red_AddRoundKeyOutput[28]), 
        .CK(clk), .Q(Red_StateRegOutput[28]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_29_ ( .D(Red_AddRoundKeyOutput[29]), 
        .CK(clk), .Q(Red_StateRegOutput[29]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_30_ ( .D(Red_AddRoundKeyOutput[30]), 
        .CK(clk), .Q(Red_StateRegOutput[30]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_31_ ( .D(Red_AddRoundKeyOutput[31]), 
        .CK(clk), .Q(Red_StateRegOutput[31]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_32_ ( .D(Red_AddRoundKeyOutput[32]), 
        .CK(clk), .Q(Red_StateRegOutput[32]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_33_ ( .D(Red_AddRoundKeyOutput[33]), 
        .CK(clk), .Q(Red_StateRegOutput[33]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_34_ ( .D(Red_AddRoundKeyOutput[34]), 
        .CK(clk), .Q(Red_StateRegOutput[34]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_35_ ( .D(Red_AddRoundKeyOutput[35]), 
        .CK(clk), .Q(Red_StateRegOutput[35]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_36_ ( .D(Red_AddRoundKeyOutput[36]), 
        .CK(clk), .Q(Red_StateRegOutput[36]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_37_ ( .D(Red_AddRoundKeyOutput[37]), 
        .CK(clk), .Q(Red_StateRegOutput[37]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_38_ ( .D(Red_AddRoundKeyOutput[38]), 
        .CK(clk), .Q(Red_StateRegOutput[38]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_39_ ( .D(Red_AddRoundKeyOutput[39]), 
        .CK(clk), .Q(Red_StateRegOutput[39]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_40_ ( .D(Red_AddRoundKeyOutput[40]), 
        .CK(clk), .Q(Red_StateRegOutput[40]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_41_ ( .D(Red_AddRoundKeyOutput[41]), 
        .CK(clk), .Q(Red_StateRegOutput[41]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_42_ ( .D(Red_AddRoundKeyOutput[42]), 
        .CK(clk), .Q(Red_StateRegOutput[42]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_43_ ( .D(Red_AddRoundKeyOutput[43]), 
        .CK(clk), .Q(Red_StateRegOutput[43]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_44_ ( .D(Red_AddRoundKeyOutput[44]), 
        .CK(clk), .Q(Red_StateRegOutput[44]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_45_ ( .D(Red_AddRoundKeyOutput[45]), 
        .CK(clk), .Q(Red_StateRegOutput[45]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_46_ ( .D(Red_AddRoundKeyOutput[46]), 
        .CK(clk), .Q(Red_StateRegOutput[46]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_47_ ( .D(Red_AddRoundKeyOutput[47]), 
        .CK(clk), .Q(Red_StateRegOutput[47]), .QN() );
  XNOR2_X1 StateRegOutputF_inst_LFInst_0_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_0_LFInst_0_n3), .B(StateRegOutput[2]), 
        .ZN(StateRegOutputF[0]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_0_LFInst_0_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[1]), .ZN(StateRegOutputF_inst_LFInst_0_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_0_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_0_LFInst_1_n3), .B(StateRegOutput[3]), 
        .ZN(StateRegOutputF[1]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_0_LFInst_1_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[1]), .ZN(StateRegOutputF_inst_LFInst_0_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_0_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_0_LFInst_2_n3), .B(StateRegOutput[3]), 
        .ZN(StateRegOutputF[2]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_0_LFInst_2_U1 ( .A(StateRegOutput[0]), 
        .B(StateRegOutput[2]), .ZN(StateRegOutputF_inst_LFInst_0_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_1_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_1_LFInst_0_n3), .B(StateRegOutput[6]), 
        .ZN(StateRegOutputF[3]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_1_LFInst_0_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[5]), .ZN(StateRegOutputF_inst_LFInst_1_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_1_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_1_LFInst_1_n3), .B(StateRegOutput[7]), 
        .ZN(StateRegOutputF[4]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_1_LFInst_1_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[5]), .ZN(StateRegOutputF_inst_LFInst_1_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_1_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_1_LFInst_2_n3), .B(StateRegOutput[7]), 
        .ZN(StateRegOutputF[5]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_1_LFInst_2_U1 ( .A(StateRegOutput[4]), 
        .B(StateRegOutput[6]), .ZN(StateRegOutputF_inst_LFInst_1_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_2_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_2_LFInst_0_n3), .B(StateRegOutput[10]), 
        .ZN(StateRegOutputF[6]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_2_LFInst_0_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[9]), .ZN(StateRegOutputF_inst_LFInst_2_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_2_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_2_LFInst_1_n3), .B(StateRegOutput[11]), 
        .ZN(StateRegOutputF[7]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_2_LFInst_1_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[9]), .ZN(StateRegOutputF_inst_LFInst_2_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_2_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_2_LFInst_2_n3), .B(StateRegOutput[11]), 
        .ZN(StateRegOutputF[8]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_2_LFInst_2_U1 ( .A(StateRegOutput[8]), 
        .B(StateRegOutput[10]), .ZN(StateRegOutputF_inst_LFInst_2_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_3_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_3_LFInst_0_n3), .B(StateRegOutput[14]), 
        .ZN(StateRegOutputF[9]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_3_LFInst_0_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[13]), .ZN(StateRegOutputF_inst_LFInst_3_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_3_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_3_LFInst_1_n3), .B(StateRegOutput[15]), 
        .ZN(StateRegOutputF[10]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_3_LFInst_1_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[13]), .ZN(StateRegOutputF_inst_LFInst_3_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_3_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_3_LFInst_2_n3), .B(StateRegOutput[15]), 
        .ZN(StateRegOutputF[11]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_3_LFInst_2_U1 ( .A(StateRegOutput[12]), 
        .B(StateRegOutput[14]), .ZN(StateRegOutputF_inst_LFInst_3_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_4_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_4_LFInst_0_n3), .B(StateRegOutput[18]), 
        .ZN(StateRegOutputF[12]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_4_LFInst_0_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[17]), .ZN(StateRegOutputF_inst_LFInst_4_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_4_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_4_LFInst_1_n3), .B(StateRegOutput[19]), 
        .ZN(StateRegOutputF[13]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_4_LFInst_1_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[17]), .ZN(StateRegOutputF_inst_LFInst_4_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_4_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_4_LFInst_2_n3), .B(StateRegOutput[19]), 
        .ZN(StateRegOutputF[14]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_4_LFInst_2_U1 ( .A(StateRegOutput[16]), 
        .B(StateRegOutput[18]), .ZN(StateRegOutputF_inst_LFInst_4_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_5_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_5_LFInst_0_n3), .B(StateRegOutput[22]), 
        .ZN(StateRegOutputF[15]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_5_LFInst_0_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[21]), .ZN(StateRegOutputF_inst_LFInst_5_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_5_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_5_LFInst_1_n3), .B(StateRegOutput[23]), 
        .ZN(StateRegOutputF[16]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_5_LFInst_1_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[21]), .ZN(StateRegOutputF_inst_LFInst_5_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_5_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_5_LFInst_2_n3), .B(StateRegOutput[23]), 
        .ZN(StateRegOutputF[17]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_5_LFInst_2_U1 ( .A(StateRegOutput[20]), 
        .B(StateRegOutput[22]), .ZN(StateRegOutputF_inst_LFInst_5_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_6_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_6_LFInst_0_n3), .B(StateRegOutput[26]), 
        .ZN(StateRegOutputF[18]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_6_LFInst_0_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[25]), .ZN(StateRegOutputF_inst_LFInst_6_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_6_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_6_LFInst_1_n3), .B(StateRegOutput[27]), 
        .ZN(StateRegOutputF[19]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_6_LFInst_1_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[25]), .ZN(StateRegOutputF_inst_LFInst_6_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_6_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_6_LFInst_2_n3), .B(StateRegOutput[27]), 
        .ZN(StateRegOutputF[20]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_6_LFInst_2_U1 ( .A(StateRegOutput[24]), 
        .B(StateRegOutput[26]), .ZN(StateRegOutputF_inst_LFInst_6_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_7_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_7_LFInst_0_n3), .B(StateRegOutput[30]), 
        .ZN(StateRegOutputF[21]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_7_LFInst_0_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[29]), .ZN(StateRegOutputF_inst_LFInst_7_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_7_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_7_LFInst_1_n3), .B(StateRegOutput[31]), 
        .ZN(StateRegOutputF[22]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_7_LFInst_1_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[29]), .ZN(StateRegOutputF_inst_LFInst_7_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_7_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_7_LFInst_2_n3), .B(StateRegOutput[31]), 
        .ZN(StateRegOutputF[23]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_7_LFInst_2_U1 ( .A(StateRegOutput[28]), 
        .B(StateRegOutput[30]), .ZN(StateRegOutputF_inst_LFInst_7_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_8_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_8_LFInst_0_n3), .B(StateRegOutput[34]), 
        .ZN(StateRegOutputF[24]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_8_LFInst_0_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[33]), .ZN(StateRegOutputF_inst_LFInst_8_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_8_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_8_LFInst_1_n3), .B(StateRegOutput[35]), 
        .ZN(StateRegOutputF[25]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_8_LFInst_1_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[33]), .ZN(StateRegOutputF_inst_LFInst_8_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_8_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_8_LFInst_2_n3), .B(StateRegOutput[35]), 
        .ZN(StateRegOutputF[26]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_8_LFInst_2_U1 ( .A(StateRegOutput[32]), 
        .B(StateRegOutput[34]), .ZN(StateRegOutputF_inst_LFInst_8_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_9_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_9_LFInst_0_n3), .B(StateRegOutput[38]), 
        .ZN(StateRegOutputF[27]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_9_LFInst_0_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[37]), .ZN(StateRegOutputF_inst_LFInst_9_LFInst_0_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_9_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_9_LFInst_1_n3), .B(StateRegOutput[39]), 
        .ZN(StateRegOutputF[28]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_9_LFInst_1_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[37]), .ZN(StateRegOutputF_inst_LFInst_9_LFInst_1_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_9_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_9_LFInst_2_n3), .B(StateRegOutput[39]), 
        .ZN(StateRegOutputF[29]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_9_LFInst_2_U1 ( .A(StateRegOutput[36]), 
        .B(StateRegOutput[38]), .ZN(StateRegOutputF_inst_LFInst_9_LFInst_2_n3)
         );
  XNOR2_X1 StateRegOutputF_inst_LFInst_10_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_10_LFInst_0_n3), .B(StateRegOutput[42]), 
        .ZN(StateRegOutputF[30]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_10_LFInst_0_U1 ( .A(StateRegOutput[40]), 
        .B(StateRegOutput[41]), .ZN(StateRegOutputF_inst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_10_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_10_LFInst_1_n3), .B(StateRegOutput[43]), 
        .ZN(StateRegOutputF[31]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_10_LFInst_1_U1 ( .A(StateRegOutput[40]), 
        .B(StateRegOutput[41]), .ZN(StateRegOutputF_inst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_10_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_10_LFInst_2_n3), .B(StateRegOutput[43]), 
        .ZN(StateRegOutputF[32]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_10_LFInst_2_U1 ( .A(StateRegOutput[40]), 
        .B(StateRegOutput[42]), .ZN(StateRegOutputF_inst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_11_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_11_LFInst_0_n3), .B(StateRegOutput[46]), 
        .ZN(StateRegOutputF[33]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_11_LFInst_0_U1 ( .A(StateRegOutput[44]), 
        .B(StateRegOutput[45]), .ZN(StateRegOutputF_inst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_11_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_11_LFInst_1_n3), .B(StateRegOutput[47]), 
        .ZN(StateRegOutputF[34]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_11_LFInst_1_U1 ( .A(StateRegOutput[44]), 
        .B(StateRegOutput[45]), .ZN(StateRegOutputF_inst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_11_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_11_LFInst_2_n3), .B(StateRegOutput[47]), 
        .ZN(StateRegOutputF[35]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_11_LFInst_2_U1 ( .A(StateRegOutput[44]), 
        .B(StateRegOutput[46]), .ZN(StateRegOutputF_inst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_12_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_12_LFInst_0_n3), .B(StateRegOutput[50]), 
        .ZN(StateRegOutputF[36]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_12_LFInst_0_U1 ( .A(StateRegOutput[48]), 
        .B(StateRegOutput[49]), .ZN(StateRegOutputF_inst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_12_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_12_LFInst_1_n3), .B(StateRegOutput[51]), 
        .ZN(StateRegOutputF[37]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_12_LFInst_1_U1 ( .A(StateRegOutput[48]), 
        .B(StateRegOutput[49]), .ZN(StateRegOutputF_inst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_12_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_12_LFInst_2_n3), .B(StateRegOutput[51]), 
        .ZN(StateRegOutputF[38]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_12_LFInst_2_U1 ( .A(StateRegOutput[48]), 
        .B(StateRegOutput[50]), .ZN(StateRegOutputF_inst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_13_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_13_LFInst_0_n3), .B(StateRegOutput[54]), 
        .ZN(StateRegOutputF[39]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_13_LFInst_0_U1 ( .A(StateRegOutput[52]), 
        .B(StateRegOutput[53]), .ZN(StateRegOutputF_inst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_13_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_13_LFInst_1_n3), .B(StateRegOutput[55]), 
        .ZN(StateRegOutputF[40]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_13_LFInst_1_U1 ( .A(StateRegOutput[52]), 
        .B(StateRegOutput[53]), .ZN(StateRegOutputF_inst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_13_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_13_LFInst_2_n3), .B(StateRegOutput[55]), 
        .ZN(StateRegOutputF[41]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_13_LFInst_2_U1 ( .A(StateRegOutput[52]), 
        .B(StateRegOutput[54]), .ZN(StateRegOutputF_inst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_14_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_14_LFInst_0_n3), .B(StateRegOutput[58]), 
        .ZN(StateRegOutputF[42]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_14_LFInst_0_U1 ( .A(StateRegOutput[56]), 
        .B(StateRegOutput[57]), .ZN(StateRegOutputF_inst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_14_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_14_LFInst_1_n3), .B(StateRegOutput[59]), 
        .ZN(StateRegOutputF[43]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_14_LFInst_1_U1 ( .A(StateRegOutput[56]), 
        .B(StateRegOutput[57]), .ZN(StateRegOutputF_inst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_14_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_14_LFInst_2_n3), .B(StateRegOutput[59]), 
        .ZN(StateRegOutputF[44]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_14_LFInst_2_U1 ( .A(StateRegOutput[56]), 
        .B(StateRegOutput[58]), .ZN(StateRegOutputF_inst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_15_LFInst_0_U2 ( .A(
        StateRegOutputF_inst_LFInst_15_LFInst_0_n3), .B(StateRegOutput[62]), 
        .ZN(StateRegOutputF[45]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_15_LFInst_0_U1 ( .A(StateRegOutput[60]), 
        .B(StateRegOutput[61]), .ZN(StateRegOutputF_inst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_15_LFInst_1_U2 ( .A(
        StateRegOutputF_inst_LFInst_15_LFInst_1_n3), .B(StateRegOutput[63]), 
        .ZN(StateRegOutputF[46]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_15_LFInst_1_U1 ( .A(StateRegOutput[60]), 
        .B(StateRegOutput[61]), .ZN(StateRegOutputF_inst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_15_LFInst_2_U2 ( .A(
        StateRegOutputF_inst_LFInst_15_LFInst_2_n3), .B(StateRegOutput[63]), 
        .ZN(StateRegOutputF[47]) );
  XNOR2_X1 StateRegOutputF_inst_LFInst_15_LFInst_2_U1 ( .A(StateRegOutput[60]), 
        .B(StateRegOutput[62]), .ZN(StateRegOutputF_inst_LFInst_15_LFInst_2_n3) );
  INV_X1 CipherErrorVecGen_XORInst_0_0_U2 ( .A(
        CipherErrorVecGen_XORInst_0_0_n6), .ZN(CipherErrorVec[0]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_0_0_U1 ( .A(StateRegOutputF[0]), .B(
        Red_StateRegOutput[0]), .ZN(CipherErrorVecGen_XORInst_0_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_0_1_U2 ( .A(
        CipherErrorVecGen_XORInst_0_1_n5), .ZN(CipherErrorVec[1]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_0_1_U1 ( .A(StateRegOutputF[1]), .B(
        Red_StateRegOutput[1]), .ZN(CipherErrorVecGen_XORInst_0_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_0_2_U2 ( .A(
        CipherErrorVecGen_XORInst_0_2_n2), .ZN(CipherErrorVec[2]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_0_2_U1 ( .A(StateRegOutputF[2]), .B(
        Red_StateRegOutput[2]), .ZN(CipherErrorVecGen_XORInst_0_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_1_0_U2 ( .A(
        CipherErrorVecGen_XORInst_1_0_n6), .ZN(CipherErrorVec[3]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_1_0_U1 ( .A(StateRegOutputF[3]), .B(
        Red_StateRegOutput[3]), .ZN(CipherErrorVecGen_XORInst_1_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_1_1_U2 ( .A(
        CipherErrorVecGen_XORInst_1_1_n5), .ZN(CipherErrorVec[4]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_1_1_U1 ( .A(StateRegOutputF[4]), .B(
        Red_StateRegOutput[4]), .ZN(CipherErrorVecGen_XORInst_1_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_1_2_U2 ( .A(
        CipherErrorVecGen_XORInst_1_2_n2), .ZN(CipherErrorVec[5]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_1_2_U1 ( .A(StateRegOutputF[5]), .B(
        Red_StateRegOutput[5]), .ZN(CipherErrorVecGen_XORInst_1_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_2_0_U2 ( .A(
        CipherErrorVecGen_XORInst_2_0_n6), .ZN(CipherErrorVec[6]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_2_0_U1 ( .A(StateRegOutputF[6]), .B(
        Red_StateRegOutput[6]), .ZN(CipherErrorVecGen_XORInst_2_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_2_1_U2 ( .A(
        CipherErrorVecGen_XORInst_2_1_n5), .ZN(CipherErrorVec[7]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_2_1_U1 ( .A(StateRegOutputF[7]), .B(
        Red_StateRegOutput[7]), .ZN(CipherErrorVecGen_XORInst_2_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_2_2_U2 ( .A(
        CipherErrorVecGen_XORInst_2_2_n2), .ZN(CipherErrorVec[8]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_2_2_U1 ( .A(StateRegOutputF[8]), .B(
        Red_StateRegOutput[8]), .ZN(CipherErrorVecGen_XORInst_2_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_3_0_U2 ( .A(
        CipherErrorVecGen_XORInst_3_0_n6), .ZN(CipherErrorVec[9]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_3_0_U1 ( .A(StateRegOutputF[9]), .B(
        Red_StateRegOutput[9]), .ZN(CipherErrorVecGen_XORInst_3_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_3_1_U2 ( .A(
        CipherErrorVecGen_XORInst_3_1_n2), .ZN(CipherErrorVec[10]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_3_1_U1 ( .A(StateRegOutputF[10]), .B(
        Red_StateRegOutput[10]), .ZN(CipherErrorVecGen_XORInst_3_1_n2) );
  INV_X1 CipherErrorVecGen_XORInst_3_2_U2 ( .A(
        CipherErrorVecGen_XORInst_3_2_n2), .ZN(CipherErrorVec[11]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_3_2_U1 ( .A(StateRegOutputF[11]), .B(
        Red_StateRegOutput[11]), .ZN(CipherErrorVecGen_XORInst_3_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_4_0_U2 ( .A(
        CipherErrorVecGen_XORInst_4_0_n6), .ZN(CipherErrorVec[12]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_4_0_U1 ( .A(StateRegOutputF[12]), .B(
        Red_StateRegOutput[12]), .ZN(CipherErrorVecGen_XORInst_4_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_4_1_U2 ( .A(
        CipherErrorVecGen_XORInst_4_1_n5), .ZN(CipherErrorVec[13]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_4_1_U1 ( .A(StateRegOutputF[13]), .B(
        Red_StateRegOutput[13]), .ZN(CipherErrorVecGen_XORInst_4_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_4_2_U2 ( .A(
        CipherErrorVecGen_XORInst_4_2_n2), .ZN(CipherErrorVec[14]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_4_2_U1 ( .A(StateRegOutputF[14]), .B(
        Red_StateRegOutput[14]), .ZN(CipherErrorVecGen_XORInst_4_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_5_0_U2 ( .A(
        CipherErrorVecGen_XORInst_5_0_n6), .ZN(CipherErrorVec[15]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_5_0_U1 ( .A(StateRegOutputF[15]), .B(
        Red_StateRegOutput[15]), .ZN(CipherErrorVecGen_XORInst_5_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_5_1_U2 ( .A(
        CipherErrorVecGen_XORInst_5_1_n5), .ZN(CipherErrorVec[16]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_5_1_U1 ( .A(StateRegOutputF[16]), .B(
        Red_StateRegOutput[16]), .ZN(CipherErrorVecGen_XORInst_5_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_5_2_U2 ( .A(
        CipherErrorVecGen_XORInst_5_2_n2), .ZN(CipherErrorVec[17]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_5_2_U1 ( .A(StateRegOutputF[17]), .B(
        Red_StateRegOutput[17]), .ZN(CipherErrorVecGen_XORInst_5_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_6_0_U2 ( .A(
        CipherErrorVecGen_XORInst_6_0_n6), .ZN(CipherErrorVec[18]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_6_0_U1 ( .A(StateRegOutputF[18]), .B(
        Red_StateRegOutput[18]), .ZN(CipherErrorVecGen_XORInst_6_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_6_1_U2 ( .A(
        CipherErrorVecGen_XORInst_6_1_n5), .ZN(CipherErrorVec[19]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_6_1_U1 ( .A(StateRegOutputF[19]), .B(
        Red_StateRegOutput[19]), .ZN(CipherErrorVecGen_XORInst_6_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_6_2_U2 ( .A(
        CipherErrorVecGen_XORInst_6_2_n2), .ZN(CipherErrorVec[20]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_6_2_U1 ( .A(StateRegOutputF[20]), .B(
        Red_StateRegOutput[20]), .ZN(CipherErrorVecGen_XORInst_6_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_7_0_U2 ( .A(
        CipherErrorVecGen_XORInst_7_0_n6), .ZN(CipherErrorVec[21]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_7_0_U1 ( .A(StateRegOutputF[21]), .B(
        Red_StateRegOutput[21]), .ZN(CipherErrorVecGen_XORInst_7_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_7_1_U2 ( .A(
        CipherErrorVecGen_XORInst_7_1_n5), .ZN(CipherErrorVec[22]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_7_1_U1 ( .A(StateRegOutputF[22]), .B(
        Red_StateRegOutput[22]), .ZN(CipherErrorVecGen_XORInst_7_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_7_2_U2 ( .A(
        CipherErrorVecGen_XORInst_7_2_n2), .ZN(CipherErrorVec[23]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_7_2_U1 ( .A(StateRegOutputF[23]), .B(
        Red_StateRegOutput[23]), .ZN(CipherErrorVecGen_XORInst_7_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_8_0_U2 ( .A(
        CipherErrorVecGen_XORInst_8_0_n6), .ZN(CipherErrorVec[24]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_8_0_U1 ( .A(StateRegOutputF[24]), .B(
        Red_StateRegOutput[24]), .ZN(CipherErrorVecGen_XORInst_8_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_8_1_U2 ( .A(
        CipherErrorVecGen_XORInst_8_1_n5), .ZN(CipherErrorVec[25]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_8_1_U1 ( .A(StateRegOutputF[25]), .B(
        Red_StateRegOutput[25]), .ZN(CipherErrorVecGen_XORInst_8_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_8_2_U2 ( .A(
        CipherErrorVecGen_XORInst_8_2_n2), .ZN(CipherErrorVec[26]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_8_2_U1 ( .A(StateRegOutputF[26]), .B(
        Red_StateRegOutput[26]), .ZN(CipherErrorVecGen_XORInst_8_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_9_0_U2 ( .A(
        CipherErrorVecGen_XORInst_9_0_n6), .ZN(CipherErrorVec[27]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_9_0_U1 ( .A(StateRegOutputF[27]), .B(
        Red_StateRegOutput[27]), .ZN(CipherErrorVecGen_XORInst_9_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_9_1_U2 ( .A(
        CipherErrorVecGen_XORInst_9_1_n5), .ZN(CipherErrorVec[28]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_9_1_U1 ( .A(StateRegOutputF[28]), .B(
        Red_StateRegOutput[28]), .ZN(CipherErrorVecGen_XORInst_9_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_9_2_U2 ( .A(
        CipherErrorVecGen_XORInst_9_2_n2), .ZN(CipherErrorVec[29]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_9_2_U1 ( .A(StateRegOutputF[29]), .B(
        Red_StateRegOutput[29]), .ZN(CipherErrorVecGen_XORInst_9_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_10_0_U2 ( .A(
        CipherErrorVecGen_XORInst_10_0_n6), .ZN(CipherErrorVec[30]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_10_0_U1 ( .A(StateRegOutputF[30]), .B(
        Red_StateRegOutput[30]), .ZN(CipherErrorVecGen_XORInst_10_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_10_1_U2 ( .A(
        CipherErrorVecGen_XORInst_10_1_n5), .ZN(CipherErrorVec[31]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_10_1_U1 ( .A(StateRegOutputF[31]), .B(
        Red_StateRegOutput[31]), .ZN(CipherErrorVecGen_XORInst_10_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_10_2_U2 ( .A(
        CipherErrorVecGen_XORInst_10_2_n2), .ZN(CipherErrorVec[32]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_10_2_U1 ( .A(StateRegOutputF[32]), .B(
        Red_StateRegOutput[32]), .ZN(CipherErrorVecGen_XORInst_10_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_11_0_U2 ( .A(
        CipherErrorVecGen_XORInst_11_0_n6), .ZN(CipherErrorVec[33]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_11_0_U1 ( .A(StateRegOutputF[33]), .B(
        Red_StateRegOutput[33]), .ZN(CipherErrorVecGen_XORInst_11_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_11_1_U2 ( .A(
        CipherErrorVecGen_XORInst_11_1_n5), .ZN(CipherErrorVec[34]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_11_1_U1 ( .A(StateRegOutputF[34]), .B(
        Red_StateRegOutput[34]), .ZN(CipherErrorVecGen_XORInst_11_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_11_2_U2 ( .A(
        CipherErrorVecGen_XORInst_11_2_n2), .ZN(CipherErrorVec[35]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_11_2_U1 ( .A(StateRegOutputF[35]), .B(
        Red_StateRegOutput[35]), .ZN(CipherErrorVecGen_XORInst_11_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_12_0_U2 ( .A(
        CipherErrorVecGen_XORInst_12_0_n6), .ZN(CipherErrorVec[36]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_12_0_U1 ( .A(StateRegOutputF[36]), .B(
        Red_StateRegOutput[36]), .ZN(CipherErrorVecGen_XORInst_12_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_12_1_U2 ( .A(
        CipherErrorVecGen_XORInst_12_1_n5), .ZN(CipherErrorVec[37]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_12_1_U1 ( .A(StateRegOutputF[37]), .B(
        Red_StateRegOutput[37]), .ZN(CipherErrorVecGen_XORInst_12_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_12_2_U2 ( .A(
        CipherErrorVecGen_XORInst_12_2_n2), .ZN(CipherErrorVec[38]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_12_2_U1 ( .A(StateRegOutputF[38]), .B(
        Red_StateRegOutput[38]), .ZN(CipherErrorVecGen_XORInst_12_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_13_0_U2 ( .A(
        CipherErrorVecGen_XORInst_13_0_n6), .ZN(CipherErrorVec[39]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_13_0_U1 ( .A(StateRegOutputF[39]), .B(
        Red_StateRegOutput[39]), .ZN(CipherErrorVecGen_XORInst_13_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_13_1_U2 ( .A(
        CipherErrorVecGen_XORInst_13_1_n5), .ZN(CipherErrorVec[40]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_13_1_U1 ( .A(StateRegOutputF[40]), .B(
        Red_StateRegOutput[40]), .ZN(CipherErrorVecGen_XORInst_13_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_13_2_U2 ( .A(
        CipherErrorVecGen_XORInst_13_2_n2), .ZN(CipherErrorVec[41]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_13_2_U1 ( .A(StateRegOutputF[41]), .B(
        Red_StateRegOutput[41]), .ZN(CipherErrorVecGen_XORInst_13_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_14_0_U2 ( .A(
        CipherErrorVecGen_XORInst_14_0_n6), .ZN(CipherErrorVec[42]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_14_0_U1 ( .A(StateRegOutputF[42]), .B(
        Red_StateRegOutput[42]), .ZN(CipherErrorVecGen_XORInst_14_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_14_1_U2 ( .A(
        CipherErrorVecGen_XORInst_14_1_n5), .ZN(CipherErrorVec[43]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_14_1_U1 ( .A(StateRegOutputF[43]), .B(
        Red_StateRegOutput[43]), .ZN(CipherErrorVecGen_XORInst_14_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_14_2_U2 ( .A(
        CipherErrorVecGen_XORInst_14_2_n2), .ZN(CipherErrorVec[44]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_14_2_U1 ( .A(StateRegOutputF[44]), .B(
        Red_StateRegOutput[44]), .ZN(CipherErrorVecGen_XORInst_14_2_n2) );
  INV_X1 CipherErrorVecGen_XORInst_15_0_U2 ( .A(
        CipherErrorVecGen_XORInst_15_0_n6), .ZN(CipherErrorVec[45]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_15_0_U1 ( .A(StateRegOutputF[45]), .B(
        Red_StateRegOutput[45]), .ZN(CipherErrorVecGen_XORInst_15_0_n6) );
  INV_X1 CipherErrorVecGen_XORInst_15_1_U2 ( .A(
        CipherErrorVecGen_XORInst_15_1_n5), .ZN(CipherErrorVec[46]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_15_1_U1 ( .A(StateRegOutputF[46]), .B(
        Red_StateRegOutput[46]), .ZN(CipherErrorVecGen_XORInst_15_1_n5) );
  INV_X1 CipherErrorVecGen_XORInst_15_2_U2 ( .A(
        CipherErrorVecGen_XORInst_15_2_n2), .ZN(CipherErrorVec[47]) );
  XNOR2_X1 CipherErrorVecGen_XORInst_15_2_U1 ( .A(StateRegOutputF[47]), .B(
        Red_StateRegOutput[47]), .ZN(CipherErrorVecGen_XORInst_15_2_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U17 ( .A(StateRegOutput[1]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n16), .ZN(Red_Feedback[45]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U15 ( .A1(CipherErrorVec[2]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U14 ( .A1(
        CipherErrorVec[1]), .A2(CipherErrorVec[0]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U11 ( .A(StateRegOutput[0]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U10 ( .A1(
        CipherErrorVec[0]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U6 ( .A(StateRegOutput[3]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U5 ( .A1(CipherErrorVec[0]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U4 ( .A1(CipherErrorVec[1]), .A2(CipherErrorVec[2]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U3 ( .A(StateRegOutput[2]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U2 ( .A1(CipherErrorVec[1]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n1), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_U1 ( .A1(CipherErrorVec[0]), .A2(CipherErrorVec[2]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_0_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n18), .ZN(Red_Feedback[46])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n10), .B(StateRegOutput[0]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U11 ( .A(CipherErrorVec[0]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U10 ( .A(StateRegOutput[2]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n7), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U9 ( .A1(CipherErrorVec[1]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U8 ( .A1(CipherErrorVec[0]), .A2(CipherErrorVec[2]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U6 ( .A(StateRegOutput[3]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U5 ( .A1(CipherErrorVec[0]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U4 ( .A1(CipherErrorVec[2]), .A2(CipherErrorVec[1]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n3), .B(StateRegOutput[1]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n2), .A2(CipherErrorVec[2]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_U1 ( .A1(CipherErrorVec[0]), .A2(CipherErrorVec[1]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_1_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n18), .ZN(Red_Feedback[47])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U17 ( .A(StateRegOutput[1]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n15), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U16 ( .A1(CipherErrorVec[2]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n7), .B(StateRegOutput[0]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U9 ( .A(CipherErrorVec[2]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U8 ( .A1(CipherErrorVec[1]), .A2(CipherErrorVec[0]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U6 ( .A(StateRegOutput[3]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U5 ( .A1(CipherErrorVec[0]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U4 ( .A1(CipherErrorVec[2]), .A2(CipherErrorVec[1]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U3 ( .A(StateRegOutput[2]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U2 ( .A1(CipherErrorVec[1]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_U1 ( .A1(CipherErrorVec[2]), .A2(CipherErrorVec[0]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_2_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U17 ( .A(StateRegOutput[5]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n16), .ZN(Red_Feedback[36]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U15 ( .A1(CipherErrorVec[5]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U14 ( .A1(
        CipherErrorVec[4]), .A2(CipherErrorVec[3]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U11 ( .A(StateRegOutput[4]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U10 ( .A1(
        CipherErrorVec[3]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U6 ( .A(StateRegOutput[7]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U5 ( .A1(CipherErrorVec[3]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U4 ( .A1(CipherErrorVec[4]), .A2(CipherErrorVec[5]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U3 ( .A(StateRegOutput[6]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U2 ( .A1(CipherErrorVec[4]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n1), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_U1 ( .A1(CipherErrorVec[3]), .A2(CipherErrorVec[5]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_3_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n18), .ZN(Red_Feedback[37])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n10), .B(StateRegOutput[4]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U11 ( .A(CipherErrorVec[3]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U10 ( .A(StateRegOutput[6]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n7), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U9 ( .A1(CipherErrorVec[4]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U8 ( .A1(CipherErrorVec[3]), .A2(CipherErrorVec[5]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U6 ( .A(StateRegOutput[7]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U5 ( .A1(CipherErrorVec[3]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U4 ( .A1(CipherErrorVec[5]), .A2(CipherErrorVec[4]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n3), .B(StateRegOutput[5]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n2), .A2(CipherErrorVec[5]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_U1 ( .A1(CipherErrorVec[3]), .A2(CipherErrorVec[4]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_4_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n18), .ZN(Red_Feedback[38])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U17 ( .A(StateRegOutput[5]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n15), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U16 ( .A1(CipherErrorVec[5]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n7), .B(StateRegOutput[4]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U9 ( .A(CipherErrorVec[5]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U8 ( .A1(CipherErrorVec[4]), .A2(CipherErrorVec[3]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U6 ( .A(StateRegOutput[7]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U5 ( .A1(CipherErrorVec[3]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U4 ( .A1(CipherErrorVec[5]), .A2(CipherErrorVec[4]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U3 ( .A(StateRegOutput[6]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U2 ( .A1(CipherErrorVec[4]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_U1 ( .A1(CipherErrorVec[5]), .A2(CipherErrorVec[3]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_5_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U17 ( .A(StateRegOutput[9]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n16), .ZN(Red_Feedback[39]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U15 ( .A1(CipherErrorVec[8]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U14 ( .A1(
        CipherErrorVec[7]), .A2(CipherErrorVec[6]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U11 ( .A(StateRegOutput[8]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U10 ( .A1(
        CipherErrorVec[6]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U6 ( .A(StateRegOutput[11]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U5 ( .A1(CipherErrorVec[6]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U4 ( .A1(CipherErrorVec[7]), .A2(CipherErrorVec[8]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U3 ( .A(StateRegOutput[10]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U2 ( .A1(CipherErrorVec[7]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n1), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_U1 ( .A1(CipherErrorVec[6]), .A2(CipherErrorVec[8]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_6_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n18), .ZN(Red_Feedback[40])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n10), .B(StateRegOutput[8]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U11 ( .A(CipherErrorVec[6]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U10 ( .A(StateRegOutput[10]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n7), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U9 ( .A1(CipherErrorVec[7]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U8 ( .A1(CipherErrorVec[6]), .A2(CipherErrorVec[8]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U6 ( .A(StateRegOutput[11]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U5 ( .A1(CipherErrorVec[6]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U4 ( .A1(CipherErrorVec[8]), .A2(CipherErrorVec[7]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n3), .B(StateRegOutput[9]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n2), .A2(CipherErrorVec[8]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_U1 ( .A1(CipherErrorVec[6]), .A2(CipherErrorVec[7]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_7_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n18), .ZN(Red_Feedback[41])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U17 ( .A(StateRegOutput[9]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n15), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U16 ( .A1(CipherErrorVec[8]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n7), .B(StateRegOutput[8]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U9 ( .A(CipherErrorVec[8]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U8 ( .A1(CipherErrorVec[7]), .A2(CipherErrorVec[6]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U6 ( .A(StateRegOutput[11]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U5 ( .A1(CipherErrorVec[6]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U4 ( .A1(CipherErrorVec[8]), .A2(CipherErrorVec[7]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U3 ( .A(StateRegOutput[10]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U2 ( .A1(CipherErrorVec[7]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_U1 ( .A1(CipherErrorVec[8]), .A2(CipherErrorVec[6]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_8_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U17 ( .A(
        StateRegOutput[13]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n16), 
        .ZN(Red_Feedback[42]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U15 ( .A1(
        CipherErrorVec[11]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n13), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U14 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U11 ( .A(
        StateRegOutput[12]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U10 ( .A1(
        CipherErrorVec[9]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U6 ( .A(StateRegOutput[15]), 
        .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U5 ( .A1(CipherErrorVec[9]), 
        .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U4 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[11]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U3 ( .A(StateRegOutput[14]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n2), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U2 ( .A1(CipherErrorVec[10]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n1), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_U1 ( .A1(CipherErrorVec[9]), .A2(CipherErrorVec[11]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_9_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n18), .ZN(Red_Feedback[43])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n10), .B(StateRegOutput[12]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U11 ( .A(CipherErrorVec[9]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U10 ( .A(
        StateRegOutput[14]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U9 ( .A1(
        CipherErrorVec[10]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U8 ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[11]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U6 ( .A(StateRegOutput[15]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U5 ( .A1(CipherErrorVec[9]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U4 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[10]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n3), .B(StateRegOutput[13]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n2), .A2(CipherErrorVec[11]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_U1 ( .A1(
        CipherErrorVec[9]), .A2(CipherErrorVec[10]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_10_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n18), .ZN(Red_Feedback[44])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U17 ( .A(
        StateRegOutput[13]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U16 ( .A1(
        CipherErrorVec[11]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n7), .B(StateRegOutput[12]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U9 ( .A(CipherErrorVec[11]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U8 ( .A1(
        CipherErrorVec[10]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U6 ( .A(StateRegOutput[15]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U5 ( .A1(CipherErrorVec[9]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U4 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[10]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U3 ( .A(StateRegOutput[14]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U2 ( .A1(
        CipherErrorVec[10]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_U1 ( .A1(
        CipherErrorVec[11]), .A2(CipherErrorVec[9]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_11_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U17 ( .A(
        StateRegOutput[17]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n16), 
        .ZN(Red_Feedback[24]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U15 ( .A1(
        CipherErrorVec[14]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U14 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U11 ( .A(
        StateRegOutput[16]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U10 ( .A1(
        CipherErrorVec[12]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U6 ( .A(StateRegOutput[19]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U5 ( .A1(
        CipherErrorVec[12]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U4 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U3 ( .A(
        StateRegOutput[18]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U2 ( .A1(
        CipherErrorVec[13]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_U1 ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_12_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n18), .ZN(Red_Feedback[25])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n10), .B(StateRegOutput[16]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U11 ( .A(CipherErrorVec[12]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U10 ( .A(
        StateRegOutput[18]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U9 ( .A1(
        CipherErrorVec[13]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U8 ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[14]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U6 ( .A(StateRegOutput[19]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U5 ( .A1(
        CipherErrorVec[12]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U4 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[13]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n3), .B(StateRegOutput[17]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n2), .A2(CipherErrorVec[14]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_U1 ( .A1(
        CipherErrorVec[12]), .A2(CipherErrorVec[13]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_13_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n18), .ZN(Red_Feedback[26])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U17 ( .A(
        StateRegOutput[17]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U16 ( .A1(
        CipherErrorVec[14]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n7), .B(StateRegOutput[16]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U9 ( .A(CipherErrorVec[14]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U8 ( .A1(
        CipherErrorVec[13]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U6 ( .A(StateRegOutput[19]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U5 ( .A1(
        CipherErrorVec[12]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U4 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[13]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U3 ( .A(StateRegOutput[18]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U2 ( .A1(
        CipherErrorVec[13]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_U1 ( .A1(
        CipherErrorVec[14]), .A2(CipherErrorVec[12]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_14_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U17 ( .A(
        StateRegOutput[21]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n16), 
        .ZN(Red_Feedback[33]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U15 ( .A1(
        CipherErrorVec[17]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U14 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U11 ( .A(
        StateRegOutput[20]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U10 ( .A1(
        CipherErrorVec[15]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U6 ( .A(StateRegOutput[23]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U5 ( .A1(
        CipherErrorVec[15]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U4 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U3 ( .A(
        StateRegOutput[22]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U2 ( .A1(
        CipherErrorVec[16]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_U1 ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_15_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n18), .ZN(Red_Feedback[34])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n10), .B(StateRegOutput[20]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U11 ( .A(CipherErrorVec[15]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U10 ( .A(
        StateRegOutput[22]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U9 ( .A1(
        CipherErrorVec[16]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U8 ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[17]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U6 ( .A(StateRegOutput[23]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U5 ( .A1(
        CipherErrorVec[15]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U4 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[16]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n3), .B(StateRegOutput[21]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n2), .A2(CipherErrorVec[17]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_U1 ( .A1(
        CipherErrorVec[15]), .A2(CipherErrorVec[16]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_16_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n18), .ZN(Red_Feedback[35])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U17 ( .A(
        StateRegOutput[21]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U16 ( .A1(
        CipherErrorVec[17]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n7), .B(StateRegOutput[20]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U9 ( .A(CipherErrorVec[17]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U8 ( .A1(
        CipherErrorVec[16]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U6 ( .A(StateRegOutput[23]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U5 ( .A1(
        CipherErrorVec[15]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U4 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[16]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U3 ( .A(StateRegOutput[22]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U2 ( .A1(
        CipherErrorVec[16]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_U1 ( .A1(
        CipherErrorVec[17]), .A2(CipherErrorVec[15]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_17_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U17 ( .A(
        StateRegOutput[25]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n16), 
        .ZN(Red_Feedback[30]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U15 ( .A1(
        CipherErrorVec[20]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U14 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U11 ( .A(
        StateRegOutput[24]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U10 ( .A1(
        CipherErrorVec[18]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U6 ( .A(StateRegOutput[27]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U5 ( .A1(
        CipherErrorVec[18]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U4 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U3 ( .A(
        StateRegOutput[26]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U2 ( .A1(
        CipherErrorVec[19]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_U1 ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_18_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n18), .ZN(Red_Feedback[31])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n10), .B(StateRegOutput[24]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U11 ( .A(CipherErrorVec[18]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U10 ( .A(
        StateRegOutput[26]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U9 ( .A1(
        CipherErrorVec[19]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U8 ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[20]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U6 ( .A(StateRegOutput[27]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U5 ( .A1(
        CipherErrorVec[18]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U4 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[19]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n3), .B(StateRegOutput[25]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n2), .A2(CipherErrorVec[20]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_U1 ( .A1(
        CipherErrorVec[18]), .A2(CipherErrorVec[19]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_19_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n18), .ZN(Red_Feedback[32])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U17 ( .A(
        StateRegOutput[25]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U16 ( .A1(
        CipherErrorVec[20]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n7), .B(StateRegOutput[24]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U9 ( .A(CipherErrorVec[20]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U8 ( .A1(
        CipherErrorVec[19]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U6 ( .A(StateRegOutput[27]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U5 ( .A1(
        CipherErrorVec[18]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U4 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[19]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U3 ( .A(StateRegOutput[26]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U2 ( .A1(
        CipherErrorVec[19]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_U1 ( .A1(
        CipherErrorVec[20]), .A2(CipherErrorVec[18]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_20_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U17 ( .A(
        StateRegOutput[29]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n16), 
        .ZN(Red_Feedback[27]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U15 ( .A1(
        CipherErrorVec[23]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U14 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U11 ( .A(
        StateRegOutput[28]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U10 ( .A1(
        CipherErrorVec[21]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U6 ( .A(StateRegOutput[31]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U5 ( .A1(
        CipherErrorVec[21]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U4 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U3 ( .A(
        StateRegOutput[30]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U2 ( .A1(
        CipherErrorVec[22]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_U1 ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_21_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n18), .ZN(Red_Feedback[28])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n10), .B(StateRegOutput[28]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U11 ( .A(CipherErrorVec[21]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U10 ( .A(
        StateRegOutput[30]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U9 ( .A1(
        CipherErrorVec[22]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U8 ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[23]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U6 ( .A(StateRegOutput[31]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U5 ( .A1(
        CipherErrorVec[21]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U4 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[22]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n3), .B(StateRegOutput[29]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n2), .A2(CipherErrorVec[23]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_U1 ( .A1(
        CipherErrorVec[21]), .A2(CipherErrorVec[22]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_22_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n18), .ZN(Red_Feedback[29])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U17 ( .A(
        StateRegOutput[29]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U16 ( .A1(
        CipherErrorVec[23]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n7), .B(StateRegOutput[28]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U9 ( .A(CipherErrorVec[23]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U8 ( .A1(
        CipherErrorVec[22]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U6 ( .A(StateRegOutput[31]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U5 ( .A1(
        CipherErrorVec[21]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U4 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[22]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U3 ( .A(StateRegOutput[30]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U2 ( .A1(
        CipherErrorVec[22]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_U1 ( .A1(
        CipherErrorVec[23]), .A2(CipherErrorVec[21]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_23_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U17 ( .A(
        StateRegOutput[33]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n16), 
        .ZN(Red_Feedback[12]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U15 ( .A1(
        CipherErrorVec[26]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U14 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U11 ( .A(
        StateRegOutput[32]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U10 ( .A1(
        CipherErrorVec[24]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U6 ( .A(StateRegOutput[35]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U5 ( .A1(
        CipherErrorVec[24]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U4 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U3 ( .A(
        StateRegOutput[34]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U2 ( .A1(
        CipherErrorVec[25]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_U1 ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_24_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n18), .ZN(Red_Feedback[13])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n10), .B(StateRegOutput[32]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U11 ( .A(CipherErrorVec[24]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U10 ( .A(
        StateRegOutput[34]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U9 ( .A1(
        CipherErrorVec[25]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U8 ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[26]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U6 ( .A(StateRegOutput[35]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U5 ( .A1(
        CipherErrorVec[24]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U4 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[25]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n3), .B(StateRegOutput[33]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n2), .A2(CipherErrorVec[26]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_U1 ( .A1(
        CipherErrorVec[24]), .A2(CipherErrorVec[25]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_25_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n18), .ZN(Red_Feedback[14])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U17 ( .A(
        StateRegOutput[33]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U16 ( .A1(
        CipherErrorVec[26]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n7), .B(StateRegOutput[32]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U9 ( .A(CipherErrorVec[26]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U8 ( .A1(
        CipherErrorVec[25]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U6 ( .A(StateRegOutput[35]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U5 ( .A1(
        CipherErrorVec[24]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U4 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[25]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U3 ( .A(StateRegOutput[34]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U2 ( .A1(
        CipherErrorVec[25]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_U1 ( .A1(
        CipherErrorVec[26]), .A2(CipherErrorVec[24]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_26_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U17 ( .A(
        StateRegOutput[37]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n16), 
        .ZN(Red_Feedback[21]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U15 ( .A1(
        CipherErrorVec[29]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U14 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U11 ( .A(
        StateRegOutput[36]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U10 ( .A1(
        CipherErrorVec[27]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U6 ( .A(StateRegOutput[39]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U5 ( .A1(
        CipherErrorVec[27]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U4 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U3 ( .A(
        StateRegOutput[38]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U2 ( .A1(
        CipherErrorVec[28]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_U1 ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_27_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n18), .ZN(Red_Feedback[22])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n10), .B(StateRegOutput[36]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U11 ( .A(CipherErrorVec[27]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U10 ( .A(
        StateRegOutput[38]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U9 ( .A1(
        CipherErrorVec[28]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U8 ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[29]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U6 ( .A(StateRegOutput[39]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U5 ( .A1(
        CipherErrorVec[27]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U4 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[28]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n3), .B(StateRegOutput[37]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n2), .A2(CipherErrorVec[29]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_U1 ( .A1(
        CipherErrorVec[27]), .A2(CipherErrorVec[28]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_28_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n18), .ZN(Red_Feedback[23])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U17 ( .A(
        StateRegOutput[37]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U16 ( .A1(
        CipherErrorVec[29]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n7), .B(StateRegOutput[36]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U9 ( .A(CipherErrorVec[29]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U8 ( .A1(
        CipherErrorVec[28]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U6 ( .A(StateRegOutput[39]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U5 ( .A1(
        CipherErrorVec[27]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U4 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[28]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U3 ( .A(StateRegOutput[38]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U2 ( .A1(
        CipherErrorVec[28]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_U1 ( .A1(
        CipherErrorVec[29]), .A2(CipherErrorVec[27]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_29_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U17 ( .A(
        StateRegOutput[41]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n16), 
        .ZN(Red_Feedback[18]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U15 ( .A1(
        CipherErrorVec[32]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U14 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U11 ( .A(
        StateRegOutput[40]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U10 ( .A1(
        CipherErrorVec[30]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U6 ( .A(StateRegOutput[43]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U5 ( .A1(
        CipherErrorVec[30]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U4 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U3 ( .A(
        StateRegOutput[42]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U2 ( .A1(
        CipherErrorVec[31]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_U1 ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_30_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n18), .ZN(Red_Feedback[19])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n10), .B(StateRegOutput[40]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U11 ( .A(CipherErrorVec[30]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U10 ( .A(
        StateRegOutput[42]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U9 ( .A1(
        CipherErrorVec[31]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U8 ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[32]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U6 ( .A(StateRegOutput[43]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U5 ( .A1(
        CipherErrorVec[30]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U4 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[31]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n3), .B(StateRegOutput[41]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n2), .A2(CipherErrorVec[32]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_U1 ( .A1(
        CipherErrorVec[30]), .A2(CipherErrorVec[31]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_31_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n18), .ZN(Red_Feedback[20])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U17 ( .A(
        StateRegOutput[41]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U16 ( .A1(
        CipherErrorVec[32]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n7), .B(StateRegOutput[40]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U9 ( .A(CipherErrorVec[32]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U8 ( .A1(
        CipherErrorVec[31]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U6 ( .A(StateRegOutput[43]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U5 ( .A1(
        CipherErrorVec[30]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U4 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[31]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U3 ( .A(StateRegOutput[42]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U2 ( .A1(
        CipherErrorVec[31]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_U1 ( .A1(
        CipherErrorVec[32]), .A2(CipherErrorVec[30]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_32_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U17 ( .A(
        StateRegOutput[45]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n16), 
        .ZN(Red_Feedback[15]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U15 ( .A1(
        CipherErrorVec[35]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U14 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U11 ( .A(
        StateRegOutput[44]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U10 ( .A1(
        CipherErrorVec[33]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U6 ( .A(StateRegOutput[47]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U5 ( .A1(
        CipherErrorVec[33]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U4 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U3 ( .A(
        StateRegOutput[46]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U2 ( .A1(
        CipherErrorVec[34]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_U1 ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_33_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n18), .ZN(Red_Feedback[16])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n10), .B(StateRegOutput[44]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U11 ( .A(CipherErrorVec[33]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U10 ( .A(
        StateRegOutput[46]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U9 ( .A1(
        CipherErrorVec[34]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U8 ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[35]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U6 ( .A(StateRegOutput[47]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U5 ( .A1(
        CipherErrorVec[33]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U4 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[34]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n3), .B(StateRegOutput[45]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n2), .A2(CipherErrorVec[35]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_U1 ( .A1(
        CipherErrorVec[33]), .A2(CipherErrorVec[34]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_34_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n18), .ZN(Red_Feedback[17])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U17 ( .A(
        StateRegOutput[45]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U16 ( .A1(
        CipherErrorVec[35]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n7), .B(StateRegOutput[44]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U9 ( .A(CipherErrorVec[35]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U8 ( .A1(
        CipherErrorVec[34]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U6 ( .A(StateRegOutput[47]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U5 ( .A1(
        CipherErrorVec[33]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U4 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[34]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U3 ( .A(StateRegOutput[46]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U2 ( .A1(
        CipherErrorVec[34]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_U1 ( .A1(
        CipherErrorVec[35]), .A2(CipherErrorVec[33]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_35_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U17 ( .A(
        StateRegOutput[49]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n16), 
        .ZN(Red_Feedback[3]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U15 ( .A1(
        CipherErrorVec[38]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U14 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U11 ( .A(
        StateRegOutput[48]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U10 ( .A1(
        CipherErrorVec[36]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U6 ( .A(StateRegOutput[51]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U5 ( .A1(
        CipherErrorVec[36]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U4 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U3 ( .A(
        StateRegOutput[50]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U2 ( .A1(
        CipherErrorVec[37]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_U1 ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_36_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n18), .ZN(Red_Feedback[4])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n10), .B(StateRegOutput[48]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U11 ( .A(CipherErrorVec[36]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U10 ( .A(
        StateRegOutput[50]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U9 ( .A1(
        CipherErrorVec[37]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U8 ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[38]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U6 ( .A(StateRegOutput[51]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U5 ( .A1(
        CipherErrorVec[36]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U4 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[37]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n3), .B(StateRegOutput[49]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n2), .A2(CipherErrorVec[38]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_U1 ( .A1(
        CipherErrorVec[36]), .A2(CipherErrorVec[37]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_37_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n18), .ZN(Red_Feedback[5])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U17 ( .A(
        StateRegOutput[49]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U16 ( .A1(
        CipherErrorVec[38]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n7), .B(StateRegOutput[48]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U9 ( .A(CipherErrorVec[38]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U8 ( .A1(
        CipherErrorVec[37]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U6 ( .A(StateRegOutput[51]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U5 ( .A1(
        CipherErrorVec[36]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U4 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[37]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U3 ( .A(StateRegOutput[50]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U2 ( .A1(
        CipherErrorVec[37]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_U1 ( .A1(
        CipherErrorVec[38]), .A2(CipherErrorVec[36]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_38_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U17 ( .A(
        StateRegOutput[53]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n16), 
        .ZN(Red_Feedback[6]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U15 ( .A1(
        CipherErrorVec[41]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U14 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U11 ( .A(
        StateRegOutput[52]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U10 ( .A1(
        CipherErrorVec[39]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U6 ( .A(StateRegOutput[55]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U5 ( .A1(
        CipherErrorVec[39]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U4 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U3 ( .A(
        StateRegOutput[54]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U2 ( .A1(
        CipherErrorVec[40]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_U1 ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_39_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n18), .ZN(Red_Feedback[7])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n10), .B(StateRegOutput[52]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U11 ( .A(CipherErrorVec[39]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U10 ( .A(
        StateRegOutput[54]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U9 ( .A1(
        CipherErrorVec[40]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U8 ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[41]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U6 ( .A(StateRegOutput[55]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U5 ( .A1(
        CipherErrorVec[39]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U4 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[40]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n3), .B(StateRegOutput[53]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n2), .A2(CipherErrorVec[41]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_U1 ( .A1(
        CipherErrorVec[39]), .A2(CipherErrorVec[40]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_40_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n18), .ZN(Red_Feedback[8])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U17 ( .A(
        StateRegOutput[53]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U16 ( .A1(
        CipherErrorVec[41]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n7), .B(StateRegOutput[52]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U9 ( .A(CipherErrorVec[41]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U8 ( .A1(
        CipherErrorVec[40]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U6 ( .A(StateRegOutput[55]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U5 ( .A1(
        CipherErrorVec[39]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U4 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[40]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U3 ( .A(StateRegOutput[54]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U2 ( .A1(
        CipherErrorVec[40]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_U1 ( .A1(
        CipherErrorVec[41]), .A2(CipherErrorVec[39]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_41_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U17 ( .A(
        StateRegOutput[57]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n16), 
        .ZN(Red_Feedback[9]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U15 ( .A1(
        CipherErrorVec[44]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U14 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U11 ( .A(
        StateRegOutput[56]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U10 ( .A1(
        CipherErrorVec[42]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U6 ( .A(StateRegOutput[59]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U5 ( .A1(
        CipherErrorVec[42]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U4 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U3 ( .A(
        StateRegOutput[58]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U2 ( .A1(
        CipherErrorVec[43]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_U1 ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_42_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n18), .ZN(Red_Feedback[10])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n10), .B(StateRegOutput[56]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U11 ( .A(CipherErrorVec[42]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U10 ( .A(
        StateRegOutput[58]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U9 ( .A1(
        CipherErrorVec[43]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U8 ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[44]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U6 ( .A(StateRegOutput[59]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U5 ( .A1(
        CipherErrorVec[42]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U4 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[43]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n3), .B(StateRegOutput[57]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n2), .A2(CipherErrorVec[44]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_U1 ( .A1(
        CipherErrorVec[42]), .A2(CipherErrorVec[43]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_43_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n18), .ZN(Red_Feedback[11])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U17 ( .A(
        StateRegOutput[57]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U16 ( .A1(
        CipherErrorVec[44]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n7), .B(StateRegOutput[56]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U9 ( .A(CipherErrorVec[44]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U8 ( .A1(
        CipherErrorVec[43]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U6 ( .A(StateRegOutput[59]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U5 ( .A1(
        CipherErrorVec[42]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U4 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[43]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U3 ( .A(StateRegOutput[58]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U2 ( .A1(
        CipherErrorVec[43]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_U1 ( .A1(
        CipherErrorVec[44]), .A2(CipherErrorVec[42]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_44_n2) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U17 ( .A(
        StateRegOutput[61]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n16), 
        .ZN(Red_Feedback[0]) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n15), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U15 ( .A1(
        CipherErrorVec[47]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n13), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n14) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U14 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n13) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U13 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n12), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n15) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n10), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U11 ( .A(
        StateRegOutput[60]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n8), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n9) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U10 ( .A1(
        CipherErrorVec[45]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n7), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n8) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U9 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U8 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n5), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n4), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U6 ( .A(StateRegOutput[63]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U5 ( .A1(
        CipherErrorVec[45]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U4 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n6) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U3 ( .A(
        StateRegOutput[62]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U2 ( .A1(
        CipherErrorVec[46]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n1), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n2) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_U1 ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_45_n1) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n18), .ZN(Red_Feedback[1])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n18) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U17 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n15), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n14), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n16) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U16 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n15) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U15 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n12), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n11), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n19) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n13), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n11) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n10), .B(StateRegOutput[60]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n9), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n8), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n10) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U11 ( .A(CipherErrorVec[45]), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U10 ( .A(
        StateRegOutput[62]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n7), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U9 ( .A1(
        CipherErrorVec[46]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n6), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n7) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U8 ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[47]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n6) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U7 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n5), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n12) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U6 ( .A(StateRegOutput[63]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n4), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n5) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U5 ( .A1(
        CipherErrorVec[45]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n9), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n4) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U4 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[46]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n9) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U3 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n3), .B(StateRegOutput[61]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n14) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U2 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n2), .A2(CipherErrorVec[47]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_U1 ( .A1(
        CipherErrorVec[45]), .A2(CipherErrorVec[46]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_46_n2) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U19 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n19), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n18), .ZN(Red_Feedback[2])
         );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U18 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n17), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n16), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n18) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U17 ( .A(
        StateRegOutput[61]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n15), 
        .Z(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n16) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U16 ( .A1(
        CipherErrorVec[47]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n14), .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n15) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U15 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n13), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n12), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n17) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U14 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n11), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n12) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U13 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n11) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U12 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n8), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n9), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n19) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U11 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n7), .B(StateRegOutput[60]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n9) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U10 ( .A1(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n14), .A2(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n6), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n7) );
  INV_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U9 ( .A(CipherErrorVec[47]), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n6) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U8 ( .A1(
        CipherErrorVec[46]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n14) );
  XNOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U7 ( .A(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n13), .B(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n10), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n8) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U6 ( .A(StateRegOutput[63]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n5), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n10) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U5 ( .A1(
        CipherErrorVec[45]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n4), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n5) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U4 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[46]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n4) );
  XOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U3 ( .A(StateRegOutput[62]), .B(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n3), .Z(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n13) );
  NOR2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U2 ( .A1(
        CipherErrorVec[46]), .A2(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n2), 
        .ZN(SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n3) );
  NAND2_X1 SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_U1 ( .A1(
        CipherErrorVec[47]), .A2(CipherErrorVec[45]), .ZN(
        SD1_Xor_FoSbox_SD1_Xor_FMulti_bit_inst_47_n2) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_0_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_0_LFInst_0_n3), .B(Feedback[2]), .ZN(
        FeedbackF[0]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_0_LFInst_0_U1 ( .A(Feedback[0]), .B(
        Feedback[1]), .ZN(StateRegOutputF_inst2_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_0_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_0_LFInst_1_n3), .B(Feedback[3]), .ZN(
        FeedbackF[1]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_0_LFInst_1_U1 ( .A(Feedback[0]), .B(
        Feedback[1]), .ZN(StateRegOutputF_inst2_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_0_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_0_LFInst_2_n3), .B(Feedback[3]), .ZN(
        FeedbackF[2]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_0_LFInst_2_U1 ( .A(Feedback[0]), .B(
        Feedback[2]), .ZN(StateRegOutputF_inst2_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_1_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_1_LFInst_0_n3), .B(Feedback[6]), .ZN(
        FeedbackF[3]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_1_LFInst_0_U1 ( .A(Feedback[4]), .B(
        Feedback[5]), .ZN(StateRegOutputF_inst2_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_1_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_1_LFInst_1_n3), .B(Feedback[7]), .ZN(
        FeedbackF[4]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_1_LFInst_1_U1 ( .A(Feedback[4]), .B(
        Feedback[5]), .ZN(StateRegOutputF_inst2_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_1_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_1_LFInst_2_n3), .B(Feedback[7]), .ZN(
        FeedbackF[5]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_1_LFInst_2_U1 ( .A(Feedback[4]), .B(
        Feedback[6]), .ZN(StateRegOutputF_inst2_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_2_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_2_LFInst_0_n3), .B(Feedback[10]), .ZN(
        FeedbackF[6]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_2_LFInst_0_U1 ( .A(Feedback[8]), .B(
        Feedback[9]), .ZN(StateRegOutputF_inst2_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_2_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_2_LFInst_1_n3), .B(Feedback[11]), .ZN(
        FeedbackF[7]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_2_LFInst_1_U1 ( .A(Feedback[8]), .B(
        Feedback[9]), .ZN(StateRegOutputF_inst2_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_2_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_2_LFInst_2_n3), .B(Feedback[11]), .ZN(
        FeedbackF[8]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_2_LFInst_2_U1 ( .A(Feedback[8]), .B(
        Feedback[10]), .ZN(StateRegOutputF_inst2_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_3_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_3_LFInst_0_n3), .B(Feedback[14]), .ZN(
        FeedbackF[9]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_3_LFInst_0_U1 ( .A(Feedback[12]), .B(
        Feedback[13]), .ZN(StateRegOutputF_inst2_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_3_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_3_LFInst_1_n3), .B(Feedback[15]), .ZN(
        FeedbackF[10]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_3_LFInst_1_U1 ( .A(Feedback[12]), .B(
        Feedback[13]), .ZN(StateRegOutputF_inst2_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_3_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_3_LFInst_2_n3), .B(Feedback[15]), .ZN(
        FeedbackF[11]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_3_LFInst_2_U1 ( .A(Feedback[12]), .B(
        Feedback[14]), .ZN(StateRegOutputF_inst2_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_4_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_4_LFInst_0_n3), .B(Feedback[18]), .ZN(
        FeedbackF[12]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_4_LFInst_0_U1 ( .A(Feedback[16]), .B(
        Feedback[17]), .ZN(StateRegOutputF_inst2_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_4_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_4_LFInst_1_n3), .B(Feedback[19]), .ZN(
        FeedbackF[13]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_4_LFInst_1_U1 ( .A(Feedback[16]), .B(
        Feedback[17]), .ZN(StateRegOutputF_inst2_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_4_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_4_LFInst_2_n3), .B(Feedback[19]), .ZN(
        FeedbackF[14]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_4_LFInst_2_U1 ( .A(Feedback[16]), .B(
        Feedback[18]), .ZN(StateRegOutputF_inst2_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_5_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_5_LFInst_0_n3), .B(Feedback[22]), .ZN(
        FeedbackF[15]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_5_LFInst_0_U1 ( .A(Feedback[20]), .B(
        Feedback[21]), .ZN(StateRegOutputF_inst2_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_5_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_5_LFInst_1_n3), .B(Feedback[23]), .ZN(
        FeedbackF[16]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_5_LFInst_1_U1 ( .A(Feedback[20]), .B(
        Feedback[21]), .ZN(StateRegOutputF_inst2_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_5_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_5_LFInst_2_n3), .B(Feedback[23]), .ZN(
        FeedbackF[17]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_5_LFInst_2_U1 ( .A(Feedback[20]), .B(
        Feedback[22]), .ZN(StateRegOutputF_inst2_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_6_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_6_LFInst_0_n3), .B(Feedback[26]), .ZN(
        FeedbackF[18]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_6_LFInst_0_U1 ( .A(Feedback[24]), .B(
        Feedback[25]), .ZN(StateRegOutputF_inst2_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_6_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_6_LFInst_1_n3), .B(Feedback[27]), .ZN(
        FeedbackF[19]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_6_LFInst_1_U1 ( .A(Feedback[24]), .B(
        Feedback[25]), .ZN(StateRegOutputF_inst2_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_6_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_6_LFInst_2_n3), .B(Feedback[27]), .ZN(
        FeedbackF[20]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_6_LFInst_2_U1 ( .A(Feedback[24]), .B(
        Feedback[26]), .ZN(StateRegOutputF_inst2_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_7_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_7_LFInst_0_n3), .B(Feedback[30]), .ZN(
        FeedbackF[21]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_7_LFInst_0_U1 ( .A(Feedback[28]), .B(
        Feedback[29]), .ZN(StateRegOutputF_inst2_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_7_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_7_LFInst_1_n3), .B(Feedback[31]), .ZN(
        FeedbackF[22]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_7_LFInst_1_U1 ( .A(Feedback[28]), .B(
        Feedback[29]), .ZN(StateRegOutputF_inst2_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_7_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_7_LFInst_2_n3), .B(Feedback[31]), .ZN(
        FeedbackF[23]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_7_LFInst_2_U1 ( .A(Feedback[28]), .B(
        Feedback[30]), .ZN(StateRegOutputF_inst2_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_8_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_8_LFInst_0_n3), .B(Feedback[34]), .ZN(
        FeedbackF[24]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_8_LFInst_0_U1 ( .A(Feedback[32]), .B(
        Feedback[33]), .ZN(StateRegOutputF_inst2_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_8_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_8_LFInst_1_n3), .B(Feedback[35]), .ZN(
        FeedbackF[25]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_8_LFInst_1_U1 ( .A(Feedback[32]), .B(
        Feedback[33]), .ZN(StateRegOutputF_inst2_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_8_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_8_LFInst_2_n3), .B(Feedback[35]), .ZN(
        FeedbackF[26]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_8_LFInst_2_U1 ( .A(Feedback[32]), .B(
        Feedback[34]), .ZN(StateRegOutputF_inst2_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_9_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_9_LFInst_0_n3), .B(Feedback[38]), .ZN(
        FeedbackF[27]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_9_LFInst_0_U1 ( .A(Feedback[36]), .B(
        Feedback[37]), .ZN(StateRegOutputF_inst2_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_9_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_9_LFInst_1_n3), .B(Feedback[39]), .ZN(
        FeedbackF[28]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_9_LFInst_1_U1 ( .A(Feedback[36]), .B(
        Feedback[37]), .ZN(StateRegOutputF_inst2_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_9_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_9_LFInst_2_n3), .B(Feedback[39]), .ZN(
        FeedbackF[29]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_9_LFInst_2_U1 ( .A(Feedback[36]), .B(
        Feedback[38]), .ZN(StateRegOutputF_inst2_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_10_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_10_LFInst_0_n3), .B(Feedback[42]), .ZN(
        FeedbackF[30]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_10_LFInst_0_U1 ( .A(Feedback[40]), .B(
        Feedback[41]), .ZN(StateRegOutputF_inst2_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_10_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_10_LFInst_1_n3), .B(Feedback[43]), .ZN(
        FeedbackF[31]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_10_LFInst_1_U1 ( .A(Feedback[40]), .B(
        Feedback[41]), .ZN(StateRegOutputF_inst2_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_10_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_10_LFInst_2_n3), .B(Feedback[43]), .ZN(
        FeedbackF[32]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_10_LFInst_2_U1 ( .A(Feedback[40]), .B(
        Feedback[42]), .ZN(StateRegOutputF_inst2_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_11_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_11_LFInst_0_n3), .B(Feedback[46]), .ZN(
        FeedbackF[33]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_11_LFInst_0_U1 ( .A(Feedback[44]), .B(
        Feedback[45]), .ZN(StateRegOutputF_inst2_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_11_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_11_LFInst_1_n3), .B(Feedback[47]), .ZN(
        FeedbackF[34]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_11_LFInst_1_U1 ( .A(Feedback[44]), .B(
        Feedback[45]), .ZN(StateRegOutputF_inst2_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_11_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_11_LFInst_2_n3), .B(Feedback[47]), .ZN(
        FeedbackF[35]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_11_LFInst_2_U1 ( .A(Feedback[44]), .B(
        Feedback[46]), .ZN(StateRegOutputF_inst2_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_12_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_12_LFInst_0_n3), .B(Feedback[50]), .ZN(
        FeedbackF[36]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_12_LFInst_0_U1 ( .A(Feedback[48]), .B(
        Feedback[49]), .ZN(StateRegOutputF_inst2_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_12_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_12_LFInst_1_n3), .B(Feedback[51]), .ZN(
        FeedbackF[37]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_12_LFInst_1_U1 ( .A(Feedback[48]), .B(
        Feedback[49]), .ZN(StateRegOutputF_inst2_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_12_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_12_LFInst_2_n3), .B(Feedback[51]), .ZN(
        FeedbackF[38]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_12_LFInst_2_U1 ( .A(Feedback[48]), .B(
        Feedback[50]), .ZN(StateRegOutputF_inst2_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_13_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_13_LFInst_0_n3), .B(Feedback[54]), .ZN(
        FeedbackF[39]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_13_LFInst_0_U1 ( .A(Feedback[52]), .B(
        Feedback[53]), .ZN(StateRegOutputF_inst2_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_13_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_13_LFInst_1_n3), .B(Feedback[55]), .ZN(
        FeedbackF[40]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_13_LFInst_1_U1 ( .A(Feedback[52]), .B(
        Feedback[53]), .ZN(StateRegOutputF_inst2_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_13_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_13_LFInst_2_n3), .B(Feedback[55]), .ZN(
        FeedbackF[41]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_13_LFInst_2_U1 ( .A(Feedback[52]), .B(
        Feedback[54]), .ZN(StateRegOutputF_inst2_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_14_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_14_LFInst_0_n3), .B(Feedback[58]), .ZN(
        FeedbackF[42]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_14_LFInst_0_U1 ( .A(Feedback[56]), .B(
        Feedback[57]), .ZN(StateRegOutputF_inst2_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_14_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_14_LFInst_1_n3), .B(Feedback[59]), .ZN(
        FeedbackF[43]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_14_LFInst_1_U1 ( .A(Feedback[56]), .B(
        Feedback[57]), .ZN(StateRegOutputF_inst2_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_14_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_14_LFInst_2_n3), .B(Feedback[59]), .ZN(
        FeedbackF[44]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_14_LFInst_2_U1 ( .A(Feedback[56]), .B(
        Feedback[58]), .ZN(StateRegOutputF_inst2_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_15_LFInst_0_U2 ( .A(
        StateRegOutputF_inst2_LFInst_15_LFInst_0_n3), .B(Feedback[62]), .ZN(
        FeedbackF[45]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_15_LFInst_0_U1 ( .A(Feedback[60]), .B(
        Feedback[61]), .ZN(StateRegOutputF_inst2_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_15_LFInst_1_U2 ( .A(
        StateRegOutputF_inst2_LFInst_15_LFInst_1_n3), .B(Feedback[63]), .ZN(
        FeedbackF[46]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_15_LFInst_1_U1 ( .A(Feedback[60]), .B(
        Feedback[61]), .ZN(StateRegOutputF_inst2_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_15_LFInst_2_U2 ( .A(
        StateRegOutputF_inst2_LFInst_15_LFInst_2_n3), .B(Feedback[63]), .ZN(
        FeedbackF[47]) );
  XNOR2_X1 StateRegOutputF_inst2_LFInst_15_LFInst_2_U1 ( .A(Feedback[60]), .B(
        Feedback[62]), .ZN(StateRegOutputF_inst2_LFInst_15_LFInst_2_n3) );
  XOR2_X1 CipherErrorVecGen2_XORInst_0_0_U1 ( .A(Red_Feedback[0]), .B(
        FeedbackF[0]), .Z(CipherErrorVec2[0]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_0_1_U1 ( .A(Red_Feedback[1]), .B(
        FeedbackF[1]), .Z(CipherErrorVec2[1]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_0_2_U1 ( .A(Red_Feedback[2]), .B(
        FeedbackF[2]), .Z(CipherErrorVec2[2]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_1_0_U1 ( .A(Red_Feedback[3]), .B(
        FeedbackF[3]), .Z(CipherErrorVec2[3]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_1_1_U1 ( .A(Red_Feedback[4]), .B(
        FeedbackF[4]), .Z(CipherErrorVec2[4]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_1_2_U1 ( .A(Red_Feedback[5]), .B(
        FeedbackF[5]), .Z(CipherErrorVec2[5]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_2_0_U1 ( .A(Red_Feedback[6]), .B(
        FeedbackF[6]), .Z(CipherErrorVec2[6]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_2_1_U1 ( .A(Red_Feedback[7]), .B(
        FeedbackF[7]), .Z(CipherErrorVec2[7]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_2_2_U1 ( .A(Red_Feedback[8]), .B(
        FeedbackF[8]), .Z(CipherErrorVec2[8]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_3_0_U1 ( .A(Red_Feedback[9]), .B(
        FeedbackF[9]), .Z(CipherErrorVec2[9]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_3_1_U1 ( .A(Red_Feedback[10]), .B(
        FeedbackF[10]), .Z(CipherErrorVec2[10]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_3_2_U1 ( .A(Red_Feedback[11]), .B(
        FeedbackF[11]), .Z(CipherErrorVec2[11]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_4_0_U1 ( .A(Red_Feedback[12]), .B(
        FeedbackF[12]), .Z(CipherErrorVec2[12]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_4_1_U1 ( .A(Red_Feedback[13]), .B(
        FeedbackF[13]), .Z(CipherErrorVec2[13]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_4_2_U1 ( .A(Red_Feedback[14]), .B(
        FeedbackF[14]), .Z(CipherErrorVec2[14]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_5_0_U1 ( .A(Red_Feedback[15]), .B(
        FeedbackF[15]), .Z(CipherErrorVec2[15]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_5_1_U1 ( .A(Red_Feedback[16]), .B(
        FeedbackF[16]), .Z(CipherErrorVec2[16]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_5_2_U1 ( .A(Red_Feedback[17]), .B(
        FeedbackF[17]), .Z(CipherErrorVec2[17]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_6_0_U1 ( .A(Red_Feedback[18]), .B(
        FeedbackF[18]), .Z(CipherErrorVec2[18]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_6_1_U1 ( .A(Red_Feedback[19]), .B(
        FeedbackF[19]), .Z(CipherErrorVec2[19]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_6_2_U1 ( .A(Red_Feedback[20]), .B(
        FeedbackF[20]), .Z(CipherErrorVec2[20]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_7_0_U1 ( .A(Red_Feedback[21]), .B(
        FeedbackF[21]), .Z(CipherErrorVec2[21]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_7_1_U1 ( .A(Red_Feedback[22]), .B(
        FeedbackF[22]), .Z(CipherErrorVec2[22]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_7_2_U1 ( .A(Red_Feedback[23]), .B(
        FeedbackF[23]), .Z(CipherErrorVec2[23]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_8_0_U1 ( .A(Red_Feedback[24]), .B(
        FeedbackF[24]), .Z(CipherErrorVec2[24]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_8_1_U1 ( .A(Red_Feedback[25]), .B(
        FeedbackF[25]), .Z(CipherErrorVec2[25]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_8_2_U1 ( .A(Red_Feedback[26]), .B(
        FeedbackF[26]), .Z(CipherErrorVec2[26]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_9_0_U1 ( .A(Red_Feedback[27]), .B(
        FeedbackF[27]), .Z(CipherErrorVec2[27]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_9_1_U1 ( .A(Red_Feedback[28]), .B(
        FeedbackF[28]), .Z(CipherErrorVec2[28]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_9_2_U1 ( .A(Red_Feedback[29]), .B(
        FeedbackF[29]), .Z(CipherErrorVec2[29]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_10_0_U1 ( .A(Red_Feedback[30]), .B(
        FeedbackF[30]), .Z(CipherErrorVec2[30]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_10_1_U1 ( .A(Red_Feedback[31]), .B(
        FeedbackF[31]), .Z(CipherErrorVec2[31]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_10_2_U1 ( .A(Red_Feedback[32]), .B(
        FeedbackF[32]), .Z(CipherErrorVec2[32]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_11_0_U1 ( .A(Red_Feedback[33]), .B(
        FeedbackF[33]), .Z(CipherErrorVec2[33]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_11_1_U1 ( .A(Red_Feedback[34]), .B(
        FeedbackF[34]), .Z(CipherErrorVec2[34]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_11_2_U1 ( .A(Red_Feedback[35]), .B(
        FeedbackF[35]), .Z(CipherErrorVec2[35]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_12_0_U1 ( .A(Red_Feedback[36]), .B(
        FeedbackF[36]), .Z(CipherErrorVec2[36]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_12_1_U1 ( .A(Red_Feedback[37]), .B(
        FeedbackF[37]), .Z(CipherErrorVec2[37]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_12_2_U1 ( .A(Red_Feedback[38]), .B(
        FeedbackF[38]), .Z(CipherErrorVec2[38]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_13_0_U1 ( .A(Red_Feedback[39]), .B(
        FeedbackF[39]), .Z(CipherErrorVec2[39]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_13_1_U1 ( .A(Red_Feedback[40]), .B(
        FeedbackF[40]), .Z(CipherErrorVec2[40]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_13_2_U1 ( .A(Red_Feedback[41]), .B(
        FeedbackF[41]), .Z(CipherErrorVec2[41]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_14_0_U1 ( .A(Red_Feedback[42]), .B(
        FeedbackF[42]), .Z(CipherErrorVec2[42]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_14_1_U1 ( .A(Red_Feedback[43]), .B(
        FeedbackF[43]), .Z(CipherErrorVec2[43]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_14_2_U1 ( .A(Red_Feedback[44]), .B(
        FeedbackF[44]), .Z(CipherErrorVec2[44]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_15_0_U1 ( .A(Red_Feedback[45]), .B(
        FeedbackF[45]), .Z(CipherErrorVec2[45]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_15_1_U1 ( .A(Red_Feedback[46]), .B(
        FeedbackF[46]), .Z(CipherErrorVec2[46]) );
  XOR2_X1 CipherErrorVecGen2_XORInst_15_2_U1 ( .A(Red_Feedback[47]), .B(
        FeedbackF[47]), .Z(CipherErrorVec2[47]) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U12 ( .A(Feedback[3]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n46), .Z(Output[3]) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U11 ( .A1(
        CipherErrorVec2[0]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U10 ( .A(Feedback[2]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n44), .ZN(Output[2])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U9 ( .A1(
        CipherErrorVec2[2]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n42), .A2(
        CipherErrorVec2[1]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U7 ( .A(Feedback[1]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n41), .ZN(Output[1])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U6 ( .A1(
        CipherErrorVec2[1]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n42), .A2(
        CipherErrorVec2[2]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U4 ( .A(Feedback[0]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n39), .Z(Output[0]) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U2 ( .A1(
        CipherErrorVec2[1]), .A2(CipherErrorVec2[2]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_U1 ( .A(
        CipherErrorVec2[0]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_0_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U12 ( .A(Feedback[7]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n46), .Z(Output[7]) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U11 ( .A1(
        CipherErrorVec2[3]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U10 ( .A(Feedback[6]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n44), .ZN(Output[6])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U9 ( .A1(
        CipherErrorVec2[5]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n42), .A2(
        CipherErrorVec2[4]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U7 ( .A(Feedback[5]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n41), .ZN(Output[5])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U6 ( .A1(
        CipherErrorVec2[4]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n42), .A2(
        CipherErrorVec2[5]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U4 ( .A(Feedback[4]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n39), .Z(Output[4]) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U2 ( .A1(
        CipherErrorVec2[4]), .A2(CipherErrorVec2[5]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_U1 ( .A(
        CipherErrorVec2[3]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_4_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U12 ( .A(Feedback[11]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n46), .Z(Output[11])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U11 ( .A1(
        CipherErrorVec2[6]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U10 ( .A(Feedback[10]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n44), .ZN(Output[10])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U9 ( .A1(
        CipherErrorVec2[8]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n42), .A2(
        CipherErrorVec2[7]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U7 ( .A(Feedback[9]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n41), .ZN(Output[9])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U6 ( .A1(
        CipherErrorVec2[7]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n42), .A2(
        CipherErrorVec2[8]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U4 ( .A(Feedback[8]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n39), .Z(Output[8]) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U2 ( .A1(
        CipherErrorVec2[7]), .A2(CipherErrorVec2[8]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_U1 ( .A(
        CipherErrorVec2[6]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_8_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U12 ( .A(Feedback[15]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n46), .Z(Output[15])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U11 ( .A1(
        CipherErrorVec2[9]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U10 ( .A(Feedback[14]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n44), .ZN(Output[14]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U9 ( .A1(
        CipherErrorVec2[11]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n42), .A2(
        CipherErrorVec2[10]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U7 ( .A(Feedback[13]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n41), .ZN(Output[13])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U6 ( .A1(
        CipherErrorVec2[10]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n42), .A2(
        CipherErrorVec2[11]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U4 ( .A(Feedback[12]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n39), .Z(Output[12])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U2 ( .A1(
        CipherErrorVec2[10]), .A2(CipherErrorVec2[11]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_U1 ( .A(
        CipherErrorVec2[9]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_12_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U12 ( .A(Feedback[19]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n46), .Z(Output[19])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U11 ( .A1(
        CipherErrorVec2[12]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U10 ( .A(Feedback[18]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n44), .ZN(Output[18]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U9 ( .A1(
        CipherErrorVec2[14]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n42), .A2(
        CipherErrorVec2[13]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U7 ( .A(Feedback[17]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n41), .ZN(Output[17])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U6 ( .A1(
        CipherErrorVec2[13]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n42), .A2(
        CipherErrorVec2[14]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U4 ( .A(Feedback[16]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n39), .Z(Output[16])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U2 ( .A1(
        CipherErrorVec2[13]), .A2(CipherErrorVec2[14]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_U1 ( .A(
        CipherErrorVec2[12]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_16_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U12 ( .A(Feedback[23]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n46), .Z(Output[23])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U11 ( .A1(
        CipherErrorVec2[15]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U10 ( .A(Feedback[22]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n44), .ZN(Output[22]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U9 ( .A1(
        CipherErrorVec2[17]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n42), .A2(
        CipherErrorVec2[16]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U7 ( .A(Feedback[21]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n41), .ZN(Output[21])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U6 ( .A1(
        CipherErrorVec2[16]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n42), .A2(
        CipherErrorVec2[17]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U4 ( .A(Feedback[20]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n39), .Z(Output[20])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U2 ( .A1(
        CipherErrorVec2[16]), .A2(CipherErrorVec2[17]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_U1 ( .A(
        CipherErrorVec2[15]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_20_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U12 ( .A(Feedback[27]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n46), .Z(Output[27])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U11 ( .A1(
        CipherErrorVec2[18]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U10 ( .A(Feedback[26]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n44), .ZN(Output[26]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U9 ( .A1(
        CipherErrorVec2[20]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n42), .A2(
        CipherErrorVec2[19]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U7 ( .A(Feedback[25]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n41), .ZN(Output[25])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U6 ( .A1(
        CipherErrorVec2[19]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n42), .A2(
        CipherErrorVec2[20]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U4 ( .A(Feedback[24]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n39), .Z(Output[24])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U2 ( .A1(
        CipherErrorVec2[19]), .A2(CipherErrorVec2[20]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_U1 ( .A(
        CipherErrorVec2[18]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_24_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U12 ( .A(Feedback[31]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n46), .Z(Output[31])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U11 ( .A1(
        CipherErrorVec2[21]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U10 ( .A(Feedback[30]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n44), .ZN(Output[30]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U9 ( .A1(
        CipherErrorVec2[23]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n42), .A2(
        CipherErrorVec2[22]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U7 ( .A(Feedback[29]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n41), .ZN(Output[29])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U6 ( .A1(
        CipherErrorVec2[22]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n42), .A2(
        CipherErrorVec2[23]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U4 ( .A(Feedback[28]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n39), .Z(Output[28])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U2 ( .A1(
        CipherErrorVec2[22]), .A2(CipherErrorVec2[23]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_U1 ( .A(
        CipherErrorVec2[21]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_28_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U12 ( .A(Feedback[35]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n46), .Z(Output[35])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U11 ( .A1(
        CipherErrorVec2[24]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U10 ( .A(Feedback[34]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n44), .ZN(Output[34]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U9 ( .A1(
        CipherErrorVec2[26]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n42), .A2(
        CipherErrorVec2[25]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U7 ( .A(Feedback[33]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n41), .ZN(Output[33])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U6 ( .A1(
        CipherErrorVec2[25]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n42), .A2(
        CipherErrorVec2[26]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U4 ( .A(Feedback[32]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n39), .Z(Output[32])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U2 ( .A1(
        CipherErrorVec2[25]), .A2(CipherErrorVec2[26]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_U1 ( .A(
        CipherErrorVec2[24]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_32_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U12 ( .A(Feedback[39]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n46), .Z(Output[39])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U11 ( .A1(
        CipherErrorVec2[27]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U10 ( .A(Feedback[38]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n44), .ZN(Output[38]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U9 ( .A1(
        CipherErrorVec2[29]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n42), .A2(
        CipherErrorVec2[28]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U7 ( .A(Feedback[37]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n41), .ZN(Output[37])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U6 ( .A1(
        CipherErrorVec2[28]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n42), .A2(
        CipherErrorVec2[29]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U4 ( .A(Feedback[36]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n39), .Z(Output[36])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U2 ( .A1(
        CipherErrorVec2[28]), .A2(CipherErrorVec2[29]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_U1 ( .A(
        CipherErrorVec2[27]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_36_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U12 ( .A(Feedback[43]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n46), .Z(Output[43])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U11 ( .A1(
        CipherErrorVec2[30]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U10 ( .A(Feedback[42]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n44), .ZN(Output[42]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U9 ( .A1(
        CipherErrorVec2[32]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n42), .A2(
        CipherErrorVec2[31]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U7 ( .A(Feedback[41]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n41), .ZN(Output[41])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U6 ( .A1(
        CipherErrorVec2[31]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n42), .A2(
        CipherErrorVec2[32]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U4 ( .A(Feedback[40]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n39), .Z(Output[40])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U2 ( .A1(
        CipherErrorVec2[31]), .A2(CipherErrorVec2[32]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_U1 ( .A(
        CipherErrorVec2[30]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_40_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U12 ( .A(Feedback[47]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n46), .Z(Output[47])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U11 ( .A1(
        CipherErrorVec2[33]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U10 ( .A(Feedback[46]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n44), .ZN(Output[46]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U9 ( .A1(
        CipherErrorVec2[35]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n42), .A2(
        CipherErrorVec2[34]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U7 ( .A(Feedback[45]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n41), .ZN(Output[45])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U6 ( .A1(
        CipherErrorVec2[34]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n42), .A2(
        CipherErrorVec2[35]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U4 ( .A(Feedback[44]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n39), .Z(Output[44])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U2 ( .A1(
        CipherErrorVec2[34]), .A2(CipherErrorVec2[35]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_U1 ( .A(
        CipherErrorVec2[33]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_44_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U12 ( .A(Feedback[51]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n46), .Z(Output[51])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U11 ( .A1(
        CipherErrorVec2[36]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U10 ( .A(Feedback[50]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n44), .ZN(Output[50]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U9 ( .A1(
        CipherErrorVec2[38]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n42), .A2(
        CipherErrorVec2[37]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U7 ( .A(Feedback[49]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n41), .ZN(Output[49])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U6 ( .A1(
        CipherErrorVec2[37]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n42), .A2(
        CipherErrorVec2[38]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U4 ( .A(Feedback[48]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n39), .Z(Output[48])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U2 ( .A1(
        CipherErrorVec2[37]), .A2(CipherErrorVec2[38]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_U1 ( .A(
        CipherErrorVec2[36]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_48_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U12 ( .A(Feedback[55]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n46), .Z(Output[55])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U11 ( .A1(
        CipherErrorVec2[39]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U10 ( .A(Feedback[54]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n44), .ZN(Output[54]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U9 ( .A1(
        CipherErrorVec2[41]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n42), .A2(
        CipherErrorVec2[40]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U7 ( .A(Feedback[53]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n41), .ZN(Output[53])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U6 ( .A1(
        CipherErrorVec2[40]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n42), .A2(
        CipherErrorVec2[41]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U4 ( .A(Feedback[52]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n39), .Z(Output[52])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U2 ( .A1(
        CipherErrorVec2[40]), .A2(CipherErrorVec2[41]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_U1 ( .A(
        CipherErrorVec2[39]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_52_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U12 ( .A(Feedback[59]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n46), .Z(Output[59])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U11 ( .A1(
        CipherErrorVec2[42]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U10 ( .A(Feedback[58]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n44), .ZN(Output[58]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U9 ( .A1(
        CipherErrorVec2[44]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n42), .A2(
        CipherErrorVec2[43]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U7 ( .A(Feedback[57]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n41), .ZN(Output[57])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U6 ( .A1(
        CipherErrorVec2[43]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n42), .A2(
        CipherErrorVec2[44]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U4 ( .A(Feedback[56]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n39), .Z(Output[56])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U2 ( .A1(
        CipherErrorVec2[43]), .A2(CipherErrorVec2[44]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_U1 ( .A(
        CipherErrorVec2[42]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_56_n42) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U12 ( .A(Feedback[63]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n46), .Z(Output[63])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U11 ( .A1(
        CipherErrorVec2[45]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n46) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U10 ( .A(Feedback[62]), .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n44), .ZN(Output[62]) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U9 ( .A1(
        CipherErrorVec2[47]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n43), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n44) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U8 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n42), .A2(
        CipherErrorVec2[46]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n43) );
  XNOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U7 ( .A(Feedback[61]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n41), .ZN(Output[61])
         );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U6 ( .A1(
        CipherErrorVec2[46]), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n40), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n41) );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U5 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n42), .A2(
        CipherErrorVec2[47]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n40) );
  XOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U4 ( .A(Feedback[60]), 
        .B(SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n39), .Z(Output[60])
         );
  NOR2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U3 ( .A1(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n42), .A2(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n45), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n39) );
  NAND2_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U2 ( .A1(
        CipherErrorVec2[46]), .A2(CipherErrorVec2[47]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n45) );
  INV_X1 SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_U1 ( .A(
        CipherErrorVec2[45]), .ZN(
        SD1_Xor_Sbox_Inst2_SD1_Xor_FMulti_bit_inst_60_n42) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_0_n3), .B(Key[2]), .ZN(Red_K1[0]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_1_n3), .B(Key[3]), .ZN(Red_K1[1]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_1_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_2_n3), .B(Key[3]), .ZN(Red_K1[2]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_2_U1 ( .A(Key[0]), .B(Key[2]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_0_n3), .B(Key[6]), .ZN(Red_K1[3]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_1_n3), .B(Key[7]), .ZN(Red_K1[4]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_1_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_2_n3), .B(Key[7]), .ZN(Red_K1[5]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_2_U1 ( .A(Key[4]), .B(Key[6]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_0_n3), .B(Key[10]), .ZN(Red_K1[6]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_1_n3), .B(Key[11]), .ZN(Red_K1[7]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_1_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_2_n3), .B(Key[11]), .ZN(Red_K1[8]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_2_U1 ( .A(Key[8]), .B(Key[10]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_0_n3), .B(Key[14]), .ZN(Red_K1[9]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_1_n3), .B(Key[15]), .ZN(Red_K1[10]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_1_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_2_n3), .B(Key[15]), .ZN(Red_K1[11]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_2_U1 ( .A(Key[12]), .B(Key[14]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_0_n3), .B(Key[18]), .ZN(Red_K1[12]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_1_n3), .B(Key[19]), .ZN(Red_K1[13]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_1_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_2_n3), .B(Key[19]), .ZN(Red_K1[14]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_2_U1 ( .A(Key[16]), .B(Key[18]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_0_n3), .B(Key[22]), .ZN(Red_K1[15]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_1_n3), .B(Key[23]), .ZN(Red_K1[16]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_1_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_2_n3), .B(Key[23]), .ZN(Red_K1[17]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_2_U1 ( .A(Key[20]), .B(Key[22]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_0_n3), .B(Key[26]), .ZN(Red_K1[18]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_1_n3), .B(Key[27]), .ZN(Red_K1[19]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_1_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_2_n3), .B(Key[27]), .ZN(Red_K1[20]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_2_U1 ( .A(Key[24]), .B(Key[26]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_0_n3), .B(Key[30]), .ZN(Red_K1[21]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_1_n3), .B(Key[31]), .ZN(Red_K1[22]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_1_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_2_n3), .B(Key[31]), .ZN(Red_K1[23]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_2_U1 ( .A(Key[28]), .B(Key[30]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_0_n3), .B(Key[34]), .ZN(Red_K1[24]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_1_n3), .B(Key[35]), .ZN(Red_K1[25]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_1_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_2_n3), .B(Key[35]), .ZN(Red_K1[26]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_2_U1 ( .A(Key[32]), .B(Key[34]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_0_n3), .B(Key[38]), .ZN(Red_K1[27]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_1_n3), .B(Key[39]), .ZN(Red_K1[28]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_1_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_2_n3), .B(Key[39]), .ZN(Red_K1[29]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_2_U1 ( .A(Key[36]), .B(Key[38]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_0_n3), .B(Key[42]), .ZN(Red_K1[30]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_1_n3), .B(Key[43]), .ZN(Red_K1[31]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_1_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_2_n3), .B(Key[43]), .ZN(Red_K1[32]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_2_U1 ( .A(Key[40]), .B(Key[42]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_0_n3), .B(Key[46]), .ZN(Red_K1[33]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_1_n3), .B(Key[47]), .ZN(Red_K1[34]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_1_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_2_n3), .B(Key[47]), .ZN(Red_K1[35]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_2_U1 ( .A(Key[44]), .B(Key[46]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_0_n3), .B(Key[50]), .ZN(Red_K1[36]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_1_n3), .B(Key[51]), .ZN(Red_K1[37]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_1_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_2_n3), .B(Key[51]), .ZN(Red_K1[38]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_2_U1 ( .A(Key[48]), .B(Key[50]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_0_n3), .B(Key[54]), .ZN(Red_K1[39]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_1_n3), .B(Key[55]), .ZN(Red_K1[40]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_1_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_2_n3), .B(Key[55]), .ZN(Red_K1[41]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_2_U1 ( .A(Key[52]), .B(Key[54]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_0_n3), .B(Key[58]), .ZN(Red_K1[42]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_1_n3), .B(Key[59]), .ZN(Red_K1[43]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_1_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_2_n3), .B(Key[59]), .ZN(Red_K1[44]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_2_U1 ( .A(Key[56]), .B(Key[58]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_0_n3), .B(Key[62]), .ZN(Red_K1[45]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_1_n3), .B(Key[63]), .ZN(Red_K1[46]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_1_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_2_n3), .B(Key[63]), .ZN(Red_K1[47]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_2_U1 ( .A(Key[60]), .B(Key[62]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_2_n3) );
endmodule

