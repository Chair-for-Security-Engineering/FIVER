
module LED64Enc ( clk, Plaintext, Key, Ciphertext, ErrorFlag );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* fiver="clock" *)input clk;
  output ErrorFlag;
  wire   Error_0_, SubCellInst_LFInst_0_LFInst_0_n7,
         SubCellInst_LFInst_0_LFInst_0_n6, SubCellInst_LFInst_0_LFInst_0_n5,
         SubCellInst_LFInst_0_LFInst_1_n26, SubCellInst_LFInst_0_LFInst_1_n25,
         SubCellInst_LFInst_0_LFInst_1_n24, SubCellInst_LFInst_0_LFInst_1_n23,
         SubCellInst_LFInst_0_LFInst_1_n22, SubCellInst_LFInst_0_LFInst_1_n21,
         SubCellInst_LFInst_0_LFInst_1_n20, SubCellInst_LFInst_0_LFInst_1_n19,
         SubCellInst_LFInst_0_LFInst_1_n18, SubCellInst_LFInst_0_LFInst_2_n28,
         SubCellInst_LFInst_0_LFInst_2_n27, SubCellInst_LFInst_0_LFInst_2_n26,
         SubCellInst_LFInst_0_LFInst_2_n25, SubCellInst_LFInst_0_LFInst_2_n24,
         SubCellInst_LFInst_0_LFInst_2_n23, SubCellInst_LFInst_0_LFInst_2_n22,
         SubCellInst_LFInst_0_LFInst_3_n26, SubCellInst_LFInst_0_LFInst_3_n25,
         SubCellInst_LFInst_0_LFInst_3_n24, SubCellInst_LFInst_0_LFInst_3_n23,
         SubCellInst_LFInst_0_LFInst_3_n22, SubCellInst_LFInst_0_LFInst_3_n21,
         SubCellInst_LFInst_0_LFInst_3_n20, SubCellInst_LFInst_0_LFInst_3_n19,
         SubCellInst_LFInst_1_LFInst_0_n7, SubCellInst_LFInst_1_LFInst_0_n6,
         SubCellInst_LFInst_1_LFInst_0_n5, SubCellInst_LFInst_1_LFInst_1_n26,
         SubCellInst_LFInst_1_LFInst_1_n25, SubCellInst_LFInst_1_LFInst_1_n24,
         SubCellInst_LFInst_1_LFInst_1_n23, SubCellInst_LFInst_1_LFInst_1_n22,
         SubCellInst_LFInst_1_LFInst_1_n21, SubCellInst_LFInst_1_LFInst_1_n20,
         SubCellInst_LFInst_1_LFInst_1_n19, SubCellInst_LFInst_1_LFInst_1_n18,
         SubCellInst_LFInst_1_LFInst_2_n28, SubCellInst_LFInst_1_LFInst_2_n27,
         SubCellInst_LFInst_1_LFInst_2_n26, SubCellInst_LFInst_1_LFInst_2_n25,
         SubCellInst_LFInst_1_LFInst_2_n24, SubCellInst_LFInst_1_LFInst_2_n23,
         SubCellInst_LFInst_1_LFInst_2_n22, SubCellInst_LFInst_1_LFInst_3_n26,
         SubCellInst_LFInst_1_LFInst_3_n25, SubCellInst_LFInst_1_LFInst_3_n24,
         SubCellInst_LFInst_1_LFInst_3_n23, SubCellInst_LFInst_1_LFInst_3_n22,
         SubCellInst_LFInst_1_LFInst_3_n21, SubCellInst_LFInst_1_LFInst_3_n20,
         SubCellInst_LFInst_1_LFInst_3_n19, SubCellInst_LFInst_2_LFInst_0_n7,
         SubCellInst_LFInst_2_LFInst_0_n6, SubCellInst_LFInst_2_LFInst_0_n5,
         SubCellInst_LFInst_2_LFInst_1_n26, SubCellInst_LFInst_2_LFInst_1_n25,
         SubCellInst_LFInst_2_LFInst_1_n24, SubCellInst_LFInst_2_LFInst_1_n23,
         SubCellInst_LFInst_2_LFInst_1_n22, SubCellInst_LFInst_2_LFInst_1_n21,
         SubCellInst_LFInst_2_LFInst_1_n20, SubCellInst_LFInst_2_LFInst_1_n19,
         SubCellInst_LFInst_2_LFInst_1_n18, SubCellInst_LFInst_2_LFInst_2_n28,
         SubCellInst_LFInst_2_LFInst_2_n27, SubCellInst_LFInst_2_LFInst_2_n26,
         SubCellInst_LFInst_2_LFInst_2_n25, SubCellInst_LFInst_2_LFInst_2_n24,
         SubCellInst_LFInst_2_LFInst_2_n23, SubCellInst_LFInst_2_LFInst_2_n22,
         SubCellInst_LFInst_2_LFInst_3_n26, SubCellInst_LFInst_2_LFInst_3_n25,
         SubCellInst_LFInst_2_LFInst_3_n24, SubCellInst_LFInst_2_LFInst_3_n23,
         SubCellInst_LFInst_2_LFInst_3_n22, SubCellInst_LFInst_2_LFInst_3_n21,
         SubCellInst_LFInst_2_LFInst_3_n20, SubCellInst_LFInst_2_LFInst_3_n19,
         SubCellInst_LFInst_3_LFInst_0_n7, SubCellInst_LFInst_3_LFInst_0_n6,
         SubCellInst_LFInst_3_LFInst_0_n5, SubCellInst_LFInst_3_LFInst_1_n26,
         SubCellInst_LFInst_3_LFInst_1_n25, SubCellInst_LFInst_3_LFInst_1_n24,
         SubCellInst_LFInst_3_LFInst_1_n23, SubCellInst_LFInst_3_LFInst_1_n22,
         SubCellInst_LFInst_3_LFInst_1_n21, SubCellInst_LFInst_3_LFInst_1_n20,
         SubCellInst_LFInst_3_LFInst_1_n19, SubCellInst_LFInst_3_LFInst_1_n18,
         SubCellInst_LFInst_3_LFInst_2_n28, SubCellInst_LFInst_3_LFInst_2_n27,
         SubCellInst_LFInst_3_LFInst_2_n26, SubCellInst_LFInst_3_LFInst_2_n25,
         SubCellInst_LFInst_3_LFInst_2_n24, SubCellInst_LFInst_3_LFInst_2_n23,
         SubCellInst_LFInst_3_LFInst_2_n22, SubCellInst_LFInst_3_LFInst_3_n26,
         SubCellInst_LFInst_3_LFInst_3_n25, SubCellInst_LFInst_3_LFInst_3_n24,
         SubCellInst_LFInst_3_LFInst_3_n23, SubCellInst_LFInst_3_LFInst_3_n22,
         SubCellInst_LFInst_3_LFInst_3_n21, SubCellInst_LFInst_3_LFInst_3_n20,
         SubCellInst_LFInst_3_LFInst_3_n19, SubCellInst_LFInst_4_LFInst_0_n7,
         SubCellInst_LFInst_4_LFInst_0_n6, SubCellInst_LFInst_4_LFInst_0_n5,
         SubCellInst_LFInst_4_LFInst_1_n26, SubCellInst_LFInst_4_LFInst_1_n25,
         SubCellInst_LFInst_4_LFInst_1_n24, SubCellInst_LFInst_4_LFInst_1_n23,
         SubCellInst_LFInst_4_LFInst_1_n22, SubCellInst_LFInst_4_LFInst_1_n21,
         SubCellInst_LFInst_4_LFInst_1_n20, SubCellInst_LFInst_4_LFInst_1_n19,
         SubCellInst_LFInst_4_LFInst_1_n18, SubCellInst_LFInst_4_LFInst_2_n28,
         SubCellInst_LFInst_4_LFInst_2_n27, SubCellInst_LFInst_4_LFInst_2_n26,
         SubCellInst_LFInst_4_LFInst_2_n25, SubCellInst_LFInst_4_LFInst_2_n24,
         SubCellInst_LFInst_4_LFInst_2_n23, SubCellInst_LFInst_4_LFInst_2_n22,
         SubCellInst_LFInst_4_LFInst_3_n26, SubCellInst_LFInst_4_LFInst_3_n25,
         SubCellInst_LFInst_4_LFInst_3_n24, SubCellInst_LFInst_4_LFInst_3_n23,
         SubCellInst_LFInst_4_LFInst_3_n22, SubCellInst_LFInst_4_LFInst_3_n21,
         SubCellInst_LFInst_4_LFInst_3_n20, SubCellInst_LFInst_4_LFInst_3_n19,
         SubCellInst_LFInst_5_LFInst_0_n7, SubCellInst_LFInst_5_LFInst_0_n6,
         SubCellInst_LFInst_5_LFInst_0_n5, SubCellInst_LFInst_5_LFInst_1_n26,
         SubCellInst_LFInst_5_LFInst_1_n25, SubCellInst_LFInst_5_LFInst_1_n24,
         SubCellInst_LFInst_5_LFInst_1_n23, SubCellInst_LFInst_5_LFInst_1_n22,
         SubCellInst_LFInst_5_LFInst_1_n21, SubCellInst_LFInst_5_LFInst_1_n20,
         SubCellInst_LFInst_5_LFInst_1_n19, SubCellInst_LFInst_5_LFInst_1_n18,
         SubCellInst_LFInst_5_LFInst_2_n28, SubCellInst_LFInst_5_LFInst_2_n27,
         SubCellInst_LFInst_5_LFInst_2_n26, SubCellInst_LFInst_5_LFInst_2_n25,
         SubCellInst_LFInst_5_LFInst_2_n24, SubCellInst_LFInst_5_LFInst_2_n23,
         SubCellInst_LFInst_5_LFInst_2_n22, SubCellInst_LFInst_5_LFInst_3_n26,
         SubCellInst_LFInst_5_LFInst_3_n25, SubCellInst_LFInst_5_LFInst_3_n24,
         SubCellInst_LFInst_5_LFInst_3_n23, SubCellInst_LFInst_5_LFInst_3_n22,
         SubCellInst_LFInst_5_LFInst_3_n21, SubCellInst_LFInst_5_LFInst_3_n20,
         SubCellInst_LFInst_5_LFInst_3_n19, SubCellInst_LFInst_6_LFInst_0_n7,
         SubCellInst_LFInst_6_LFInst_0_n6, SubCellInst_LFInst_6_LFInst_0_n5,
         SubCellInst_LFInst_6_LFInst_1_n26, SubCellInst_LFInst_6_LFInst_1_n25,
         SubCellInst_LFInst_6_LFInst_1_n24, SubCellInst_LFInst_6_LFInst_1_n23,
         SubCellInst_LFInst_6_LFInst_1_n22, SubCellInst_LFInst_6_LFInst_1_n21,
         SubCellInst_LFInst_6_LFInst_1_n20, SubCellInst_LFInst_6_LFInst_1_n19,
         SubCellInst_LFInst_6_LFInst_1_n18, SubCellInst_LFInst_6_LFInst_2_n28,
         SubCellInst_LFInst_6_LFInst_2_n27, SubCellInst_LFInst_6_LFInst_2_n26,
         SubCellInst_LFInst_6_LFInst_2_n25, SubCellInst_LFInst_6_LFInst_2_n24,
         SubCellInst_LFInst_6_LFInst_2_n23, SubCellInst_LFInst_6_LFInst_2_n22,
         SubCellInst_LFInst_6_LFInst_3_n26, SubCellInst_LFInst_6_LFInst_3_n25,
         SubCellInst_LFInst_6_LFInst_3_n24, SubCellInst_LFInst_6_LFInst_3_n23,
         SubCellInst_LFInst_6_LFInst_3_n22, SubCellInst_LFInst_6_LFInst_3_n21,
         SubCellInst_LFInst_6_LFInst_3_n20, SubCellInst_LFInst_6_LFInst_3_n19,
         SubCellInst_LFInst_7_LFInst_0_n7, SubCellInst_LFInst_7_LFInst_0_n6,
         SubCellInst_LFInst_7_LFInst_0_n5, SubCellInst_LFInst_7_LFInst_1_n26,
         SubCellInst_LFInst_7_LFInst_1_n25, SubCellInst_LFInst_7_LFInst_1_n24,
         SubCellInst_LFInst_7_LFInst_1_n23, SubCellInst_LFInst_7_LFInst_1_n22,
         SubCellInst_LFInst_7_LFInst_1_n21, SubCellInst_LFInst_7_LFInst_1_n20,
         SubCellInst_LFInst_7_LFInst_1_n19, SubCellInst_LFInst_7_LFInst_1_n18,
         SubCellInst_LFInst_7_LFInst_2_n28, SubCellInst_LFInst_7_LFInst_2_n27,
         SubCellInst_LFInst_7_LFInst_2_n26, SubCellInst_LFInst_7_LFInst_2_n25,
         SubCellInst_LFInst_7_LFInst_2_n24, SubCellInst_LFInst_7_LFInst_2_n23,
         SubCellInst_LFInst_7_LFInst_2_n22, SubCellInst_LFInst_7_LFInst_3_n26,
         SubCellInst_LFInst_7_LFInst_3_n25, SubCellInst_LFInst_7_LFInst_3_n24,
         SubCellInst_LFInst_7_LFInst_3_n23, SubCellInst_LFInst_7_LFInst_3_n22,
         SubCellInst_LFInst_7_LFInst_3_n21, SubCellInst_LFInst_7_LFInst_3_n20,
         SubCellInst_LFInst_7_LFInst_3_n19, SubCellInst_LFInst_8_LFInst_0_n7,
         SubCellInst_LFInst_8_LFInst_0_n6, SubCellInst_LFInst_8_LFInst_0_n5,
         SubCellInst_LFInst_8_LFInst_1_n26, SubCellInst_LFInst_8_LFInst_1_n25,
         SubCellInst_LFInst_8_LFInst_1_n24, SubCellInst_LFInst_8_LFInst_1_n23,
         SubCellInst_LFInst_8_LFInst_1_n22, SubCellInst_LFInst_8_LFInst_1_n21,
         SubCellInst_LFInst_8_LFInst_1_n20, SubCellInst_LFInst_8_LFInst_1_n19,
         SubCellInst_LFInst_8_LFInst_1_n18, SubCellInst_LFInst_8_LFInst_2_n28,
         SubCellInst_LFInst_8_LFInst_2_n27, SubCellInst_LFInst_8_LFInst_2_n26,
         SubCellInst_LFInst_8_LFInst_2_n25, SubCellInst_LFInst_8_LFInst_2_n24,
         SubCellInst_LFInst_8_LFInst_2_n23, SubCellInst_LFInst_8_LFInst_2_n22,
         SubCellInst_LFInst_8_LFInst_3_n26, SubCellInst_LFInst_8_LFInst_3_n25,
         SubCellInst_LFInst_8_LFInst_3_n24, SubCellInst_LFInst_8_LFInst_3_n23,
         SubCellInst_LFInst_8_LFInst_3_n22, SubCellInst_LFInst_8_LFInst_3_n21,
         SubCellInst_LFInst_8_LFInst_3_n20, SubCellInst_LFInst_8_LFInst_3_n19,
         SubCellInst_LFInst_9_LFInst_0_n7, SubCellInst_LFInst_9_LFInst_0_n6,
         SubCellInst_LFInst_9_LFInst_0_n5, SubCellInst_LFInst_9_LFInst_1_n26,
         SubCellInst_LFInst_9_LFInst_1_n25, SubCellInst_LFInst_9_LFInst_1_n24,
         SubCellInst_LFInst_9_LFInst_1_n23, SubCellInst_LFInst_9_LFInst_1_n22,
         SubCellInst_LFInst_9_LFInst_1_n21, SubCellInst_LFInst_9_LFInst_1_n20,
         SubCellInst_LFInst_9_LFInst_1_n19, SubCellInst_LFInst_9_LFInst_1_n18,
         SubCellInst_LFInst_9_LFInst_2_n28, SubCellInst_LFInst_9_LFInst_2_n27,
         SubCellInst_LFInst_9_LFInst_2_n26, SubCellInst_LFInst_9_LFInst_2_n25,
         SubCellInst_LFInst_9_LFInst_2_n24, SubCellInst_LFInst_9_LFInst_2_n23,
         SubCellInst_LFInst_9_LFInst_2_n22, SubCellInst_LFInst_9_LFInst_3_n26,
         SubCellInst_LFInst_9_LFInst_3_n25, SubCellInst_LFInst_9_LFInst_3_n24,
         SubCellInst_LFInst_9_LFInst_3_n23, SubCellInst_LFInst_9_LFInst_3_n22,
         SubCellInst_LFInst_9_LFInst_3_n21, SubCellInst_LFInst_9_LFInst_3_n20,
         SubCellInst_LFInst_9_LFInst_3_n19, SubCellInst_LFInst_10_LFInst_0_n7,
         SubCellInst_LFInst_10_LFInst_0_n6, SubCellInst_LFInst_10_LFInst_0_n5,
         SubCellInst_LFInst_10_LFInst_1_n26,
         SubCellInst_LFInst_10_LFInst_1_n25,
         SubCellInst_LFInst_10_LFInst_1_n24,
         SubCellInst_LFInst_10_LFInst_1_n23,
         SubCellInst_LFInst_10_LFInst_1_n22,
         SubCellInst_LFInst_10_LFInst_1_n21,
         SubCellInst_LFInst_10_LFInst_1_n20,
         SubCellInst_LFInst_10_LFInst_1_n19,
         SubCellInst_LFInst_10_LFInst_1_n18,
         SubCellInst_LFInst_10_LFInst_2_n28,
         SubCellInst_LFInst_10_LFInst_2_n27,
         SubCellInst_LFInst_10_LFInst_2_n26,
         SubCellInst_LFInst_10_LFInst_2_n25,
         SubCellInst_LFInst_10_LFInst_2_n24,
         SubCellInst_LFInst_10_LFInst_2_n23,
         SubCellInst_LFInst_10_LFInst_2_n22,
         SubCellInst_LFInst_10_LFInst_3_n26,
         SubCellInst_LFInst_10_LFInst_3_n25,
         SubCellInst_LFInst_10_LFInst_3_n24,
         SubCellInst_LFInst_10_LFInst_3_n23,
         SubCellInst_LFInst_10_LFInst_3_n22,
         SubCellInst_LFInst_10_LFInst_3_n21,
         SubCellInst_LFInst_10_LFInst_3_n20,
         SubCellInst_LFInst_10_LFInst_3_n19, SubCellInst_LFInst_11_LFInst_0_n7,
         SubCellInst_LFInst_11_LFInst_0_n6, SubCellInst_LFInst_11_LFInst_0_n5,
         SubCellInst_LFInst_11_LFInst_1_n26,
         SubCellInst_LFInst_11_LFInst_1_n25,
         SubCellInst_LFInst_11_LFInst_1_n24,
         SubCellInst_LFInst_11_LFInst_1_n23,
         SubCellInst_LFInst_11_LFInst_1_n22,
         SubCellInst_LFInst_11_LFInst_1_n21,
         SubCellInst_LFInst_11_LFInst_1_n20,
         SubCellInst_LFInst_11_LFInst_1_n19,
         SubCellInst_LFInst_11_LFInst_1_n18,
         SubCellInst_LFInst_11_LFInst_2_n28,
         SubCellInst_LFInst_11_LFInst_2_n27,
         SubCellInst_LFInst_11_LFInst_2_n26,
         SubCellInst_LFInst_11_LFInst_2_n25,
         SubCellInst_LFInst_11_LFInst_2_n24,
         SubCellInst_LFInst_11_LFInst_2_n23,
         SubCellInst_LFInst_11_LFInst_2_n22,
         SubCellInst_LFInst_11_LFInst_3_n26,
         SubCellInst_LFInst_11_LFInst_3_n25,
         SubCellInst_LFInst_11_LFInst_3_n24,
         SubCellInst_LFInst_11_LFInst_3_n23,
         SubCellInst_LFInst_11_LFInst_3_n22,
         SubCellInst_LFInst_11_LFInst_3_n21,
         SubCellInst_LFInst_11_LFInst_3_n20,
         SubCellInst_LFInst_11_LFInst_3_n19, SubCellInst_LFInst_12_LFInst_0_n7,
         SubCellInst_LFInst_12_LFInst_0_n6, SubCellInst_LFInst_12_LFInst_0_n5,
         SubCellInst_LFInst_12_LFInst_1_n26,
         SubCellInst_LFInst_12_LFInst_1_n25,
         SubCellInst_LFInst_12_LFInst_1_n24,
         SubCellInst_LFInst_12_LFInst_1_n23,
         SubCellInst_LFInst_12_LFInst_1_n22,
         SubCellInst_LFInst_12_LFInst_1_n21,
         SubCellInst_LFInst_12_LFInst_1_n20,
         SubCellInst_LFInst_12_LFInst_1_n19,
         SubCellInst_LFInst_12_LFInst_1_n18,
         SubCellInst_LFInst_12_LFInst_2_n28,
         SubCellInst_LFInst_12_LFInst_2_n27,
         SubCellInst_LFInst_12_LFInst_2_n26,
         SubCellInst_LFInst_12_LFInst_2_n25,
         SubCellInst_LFInst_12_LFInst_2_n24,
         SubCellInst_LFInst_12_LFInst_2_n23,
         SubCellInst_LFInst_12_LFInst_2_n22,
         SubCellInst_LFInst_12_LFInst_3_n26,
         SubCellInst_LFInst_12_LFInst_3_n25,
         SubCellInst_LFInst_12_LFInst_3_n24,
         SubCellInst_LFInst_12_LFInst_3_n23,
         SubCellInst_LFInst_12_LFInst_3_n22,
         SubCellInst_LFInst_12_LFInst_3_n21,
         SubCellInst_LFInst_12_LFInst_3_n20,
         SubCellInst_LFInst_12_LFInst_3_n19, SubCellInst_LFInst_13_LFInst_0_n7,
         SubCellInst_LFInst_13_LFInst_0_n6, SubCellInst_LFInst_13_LFInst_0_n5,
         SubCellInst_LFInst_13_LFInst_1_n26,
         SubCellInst_LFInst_13_LFInst_1_n25,
         SubCellInst_LFInst_13_LFInst_1_n24,
         SubCellInst_LFInst_13_LFInst_1_n23,
         SubCellInst_LFInst_13_LFInst_1_n22,
         SubCellInst_LFInst_13_LFInst_1_n21,
         SubCellInst_LFInst_13_LFInst_1_n20,
         SubCellInst_LFInst_13_LFInst_1_n19,
         SubCellInst_LFInst_13_LFInst_1_n18,
         SubCellInst_LFInst_13_LFInst_2_n28,
         SubCellInst_LFInst_13_LFInst_2_n27,
         SubCellInst_LFInst_13_LFInst_2_n26,
         SubCellInst_LFInst_13_LFInst_2_n25,
         SubCellInst_LFInst_13_LFInst_2_n24,
         SubCellInst_LFInst_13_LFInst_2_n23,
         SubCellInst_LFInst_13_LFInst_2_n22,
         SubCellInst_LFInst_13_LFInst_3_n26,
         SubCellInst_LFInst_13_LFInst_3_n25,
         SubCellInst_LFInst_13_LFInst_3_n24,
         SubCellInst_LFInst_13_LFInst_3_n23,
         SubCellInst_LFInst_13_LFInst_3_n22,
         SubCellInst_LFInst_13_LFInst_3_n21,
         SubCellInst_LFInst_13_LFInst_3_n20,
         SubCellInst_LFInst_13_LFInst_3_n19, SubCellInst_LFInst_14_LFInst_0_n7,
         SubCellInst_LFInst_14_LFInst_0_n6, SubCellInst_LFInst_14_LFInst_0_n5,
         SubCellInst_LFInst_14_LFInst_1_n26,
         SubCellInst_LFInst_14_LFInst_1_n25,
         SubCellInst_LFInst_14_LFInst_1_n24,
         SubCellInst_LFInst_14_LFInst_1_n23,
         SubCellInst_LFInst_14_LFInst_1_n22,
         SubCellInst_LFInst_14_LFInst_1_n21,
         SubCellInst_LFInst_14_LFInst_1_n20,
         SubCellInst_LFInst_14_LFInst_1_n19,
         SubCellInst_LFInst_14_LFInst_1_n18,
         SubCellInst_LFInst_14_LFInst_2_n28,
         SubCellInst_LFInst_14_LFInst_2_n27,
         SubCellInst_LFInst_14_LFInst_2_n26,
         SubCellInst_LFInst_14_LFInst_2_n25,
         SubCellInst_LFInst_14_LFInst_2_n24,
         SubCellInst_LFInst_14_LFInst_2_n23,
         SubCellInst_LFInst_14_LFInst_2_n22,
         SubCellInst_LFInst_14_LFInst_3_n26,
         SubCellInst_LFInst_14_LFInst_3_n25,
         SubCellInst_LFInst_14_LFInst_3_n24,
         SubCellInst_LFInst_14_LFInst_3_n23,
         SubCellInst_LFInst_14_LFInst_3_n22,
         SubCellInst_LFInst_14_LFInst_3_n21,
         SubCellInst_LFInst_14_LFInst_3_n20,
         SubCellInst_LFInst_14_LFInst_3_n19, SubCellInst_LFInst_15_LFInst_0_n7,
         SubCellInst_LFInst_15_LFInst_0_n6, SubCellInst_LFInst_15_LFInst_0_n5,
         SubCellInst_LFInst_15_LFInst_1_n26,
         SubCellInst_LFInst_15_LFInst_1_n25,
         SubCellInst_LFInst_15_LFInst_1_n24,
         SubCellInst_LFInst_15_LFInst_1_n23,
         SubCellInst_LFInst_15_LFInst_1_n22,
         SubCellInst_LFInst_15_LFInst_1_n21,
         SubCellInst_LFInst_15_LFInst_1_n20,
         SubCellInst_LFInst_15_LFInst_1_n19,
         SubCellInst_LFInst_15_LFInst_1_n18,
         SubCellInst_LFInst_15_LFInst_2_n28,
         SubCellInst_LFInst_15_LFInst_2_n27,
         SubCellInst_LFInst_15_LFInst_2_n26,
         SubCellInst_LFInst_15_LFInst_2_n25,
         SubCellInst_LFInst_15_LFInst_2_n24,
         SubCellInst_LFInst_15_LFInst_2_n23,
         SubCellInst_LFInst_15_LFInst_2_n22,
         SubCellInst_LFInst_15_LFInst_3_n26,
         SubCellInst_LFInst_15_LFInst_3_n25,
         SubCellInst_LFInst_15_LFInst_3_n24,
         SubCellInst_LFInst_15_LFInst_3_n23,
         SubCellInst_LFInst_15_LFInst_3_n22,
         SubCellInst_LFInst_15_LFInst_3_n21,
         SubCellInst_LFInst_15_LFInst_3_n20,
         SubCellInst_LFInst_15_LFInst_3_n19, MCInst_MC0_v0_2Inst_0_n3,
         MCInst_MC0_v1_2Inst_0_n3, MCInst_MC0_v2_3Inst_0_n6,
         MCInst_MC0_v2_3Inst_0_n5, MCInst_MC0_v3_3Inst_0_n3,
         MCInst_MC0_v0_2Inst_1_n3, MCInst_MC0_v2_1Inst_1_n3,
         MCInst_MC0_v2_2Inst_1_n6, MCInst_MC0_v2_2Inst_1_n5,
         MCInst_MC0_v3_3Inst_1_n3, MCInst_MC0_v1_1Inst_2_n3,
         MCInst_MC0_v1_2Inst_2_n3, MCInst_MC0_v2_1Inst_2_n3,
         MCInst_MC0_v2_2Inst_2_n3, MCInst_MC0_v3_1Inst_2_n3,
         MCInst_MC0_v1_2Inst_3_n6, MCInst_MC0_v1_2Inst_3_n5,
         MCInst_MC0_v2_2Inst_3_n3, MCInst_MC0_v2_3Inst_3_n3,
         MCInst_MC0_r0Inst_XORInst_0_0_n8, MCInst_MC0_r0Inst_XORInst_0_0_n7,
         MCInst_MC0_r0Inst_XORInst_0_1_n8, MCInst_MC0_r0Inst_XORInst_0_1_n7,
         MCInst_MC0_r0Inst_XORInst_0_2_n8, MCInst_MC0_r0Inst_XORInst_0_2_n7,
         MCInst_MC0_r0Inst_XORInst_0_3_n8, MCInst_MC0_r0Inst_XORInst_0_3_n7,
         MCInst_MC0_r1Inst_XORInst_0_0_n8, MCInst_MC0_r1Inst_XORInst_0_0_n7,
         MCInst_MC0_r1Inst_XORInst_0_1_n8, MCInst_MC0_r1Inst_XORInst_0_1_n7,
         MCInst_MC0_r1Inst_XORInst_0_2_n8, MCInst_MC0_r1Inst_XORInst_0_2_n7,
         MCInst_MC0_r1Inst_XORInst_0_3_n8, MCInst_MC0_r1Inst_XORInst_0_3_n7,
         MCInst_MC0_r2Inst_XORInst_0_0_n8, MCInst_MC0_r2Inst_XORInst_0_0_n7,
         MCInst_MC0_r2Inst_XORInst_0_1_n8, MCInst_MC0_r2Inst_XORInst_0_1_n7,
         MCInst_MC0_r2Inst_XORInst_0_2_n8, MCInst_MC0_r2Inst_XORInst_0_2_n7,
         MCInst_MC0_r2Inst_XORInst_0_3_n8, MCInst_MC0_r2Inst_XORInst_0_3_n7,
         MCInst_MC0_r3Inst_XORInst_0_0_n8, MCInst_MC0_r3Inst_XORInst_0_0_n7,
         MCInst_MC0_r3Inst_XORInst_0_1_n8, MCInst_MC0_r3Inst_XORInst_0_1_n7,
         MCInst_MC0_r3Inst_XORInst_0_2_n8, MCInst_MC0_r3Inst_XORInst_0_2_n7,
         MCInst_MC0_r3Inst_XORInst_0_3_n8, MCInst_MC0_r3Inst_XORInst_0_3_n7,
         MCInst_MC1_v0_2Inst_0_n3, MCInst_MC1_v1_2Inst_0_n3,
         MCInst_MC1_v2_3Inst_0_n6, MCInst_MC1_v2_3Inst_0_n5,
         MCInst_MC1_v3_3Inst_0_n3, MCInst_MC1_v0_2Inst_1_n3,
         MCInst_MC1_v2_1Inst_1_n3, MCInst_MC1_v2_2Inst_1_n6,
         MCInst_MC1_v2_2Inst_1_n5, MCInst_MC1_v3_3Inst_1_n3,
         MCInst_MC1_v1_1Inst_2_n3, MCInst_MC1_v1_2Inst_2_n3,
         MCInst_MC1_v2_1Inst_2_n3, MCInst_MC1_v2_2Inst_2_n3,
         MCInst_MC1_v3_1Inst_2_n3, MCInst_MC1_v1_2Inst_3_n6,
         MCInst_MC1_v1_2Inst_3_n5, MCInst_MC1_v2_2Inst_3_n3,
         MCInst_MC1_v2_3Inst_3_n3, MCInst_MC1_r0Inst_XORInst_0_0_n8,
         MCInst_MC1_r0Inst_XORInst_0_0_n7, MCInst_MC1_r0Inst_XORInst_0_1_n8,
         MCInst_MC1_r0Inst_XORInst_0_1_n7, MCInst_MC1_r0Inst_XORInst_0_2_n8,
         MCInst_MC1_r0Inst_XORInst_0_2_n7, MCInst_MC1_r0Inst_XORInst_0_3_n8,
         MCInst_MC1_r0Inst_XORInst_0_3_n7, MCInst_MC1_r1Inst_XORInst_0_0_n8,
         MCInst_MC1_r1Inst_XORInst_0_0_n7, MCInst_MC1_r1Inst_XORInst_0_1_n8,
         MCInst_MC1_r1Inst_XORInst_0_1_n7, MCInst_MC1_r1Inst_XORInst_0_2_n8,
         MCInst_MC1_r1Inst_XORInst_0_2_n7, MCInst_MC1_r1Inst_XORInst_0_3_n8,
         MCInst_MC1_r1Inst_XORInst_0_3_n7, MCInst_MC1_r2Inst_XORInst_0_0_n8,
         MCInst_MC1_r2Inst_XORInst_0_0_n7, MCInst_MC1_r2Inst_XORInst_0_1_n8,
         MCInst_MC1_r2Inst_XORInst_0_1_n7, MCInst_MC1_r2Inst_XORInst_0_2_n8,
         MCInst_MC1_r2Inst_XORInst_0_2_n7, MCInst_MC1_r2Inst_XORInst_0_3_n8,
         MCInst_MC1_r2Inst_XORInst_0_3_n7, MCInst_MC1_r3Inst_XORInst_0_0_n8,
         MCInst_MC1_r3Inst_XORInst_0_0_n7, MCInst_MC1_r3Inst_XORInst_0_1_n8,
         MCInst_MC1_r3Inst_XORInst_0_1_n7, MCInst_MC1_r3Inst_XORInst_0_2_n8,
         MCInst_MC1_r3Inst_XORInst_0_2_n7, MCInst_MC1_r3Inst_XORInst_0_3_n8,
         MCInst_MC1_r3Inst_XORInst_0_3_n7, MCInst_MC2_v0_2Inst_0_n3,
         MCInst_MC2_v1_2Inst_0_n3, MCInst_MC2_v2_3Inst_0_n6,
         MCInst_MC2_v2_3Inst_0_n5, MCInst_MC2_v3_3Inst_0_n3,
         MCInst_MC2_v0_2Inst_1_n3, MCInst_MC2_v2_1Inst_1_n3,
         MCInst_MC2_v2_2Inst_1_n6, MCInst_MC2_v2_2Inst_1_n5,
         MCInst_MC2_v3_3Inst_1_n3, MCInst_MC2_v1_1Inst_2_n3,
         MCInst_MC2_v1_2Inst_2_n3, MCInst_MC2_v2_1Inst_2_n3,
         MCInst_MC2_v2_2Inst_2_n3, MCInst_MC2_v3_1Inst_2_n3,
         MCInst_MC2_v1_2Inst_3_n6, MCInst_MC2_v1_2Inst_3_n5,
         MCInst_MC2_v2_2Inst_3_n3, MCInst_MC2_v2_3Inst_3_n3,
         MCInst_MC2_r0Inst_XORInst_0_0_n8, MCInst_MC2_r0Inst_XORInst_0_0_n7,
         MCInst_MC2_r0Inst_XORInst_0_1_n8, MCInst_MC2_r0Inst_XORInst_0_1_n7,
         MCInst_MC2_r0Inst_XORInst_0_2_n8, MCInst_MC2_r0Inst_XORInst_0_2_n7,
         MCInst_MC2_r0Inst_XORInst_0_3_n8, MCInst_MC2_r0Inst_XORInst_0_3_n7,
         MCInst_MC2_r1Inst_XORInst_0_0_n8, MCInst_MC2_r1Inst_XORInst_0_0_n7,
         MCInst_MC2_r1Inst_XORInst_0_1_n8, MCInst_MC2_r1Inst_XORInst_0_1_n7,
         MCInst_MC2_r1Inst_XORInst_0_2_n8, MCInst_MC2_r1Inst_XORInst_0_2_n7,
         MCInst_MC2_r1Inst_XORInst_0_3_n8, MCInst_MC2_r1Inst_XORInst_0_3_n7,
         MCInst_MC2_r2Inst_XORInst_0_0_n8, MCInst_MC2_r2Inst_XORInst_0_0_n7,
         MCInst_MC2_r2Inst_XORInst_0_1_n8, MCInst_MC2_r2Inst_XORInst_0_1_n7,
         MCInst_MC2_r2Inst_XORInst_0_2_n8, MCInst_MC2_r2Inst_XORInst_0_2_n7,
         MCInst_MC2_r2Inst_XORInst_0_3_n8, MCInst_MC2_r2Inst_XORInst_0_3_n7,
         MCInst_MC2_r3Inst_XORInst_0_0_n8, MCInst_MC2_r3Inst_XORInst_0_0_n7,
         MCInst_MC2_r3Inst_XORInst_0_1_n8, MCInst_MC2_r3Inst_XORInst_0_1_n7,
         MCInst_MC2_r3Inst_XORInst_0_2_n8, MCInst_MC2_r3Inst_XORInst_0_2_n7,
         MCInst_MC2_r3Inst_XORInst_0_3_n8, MCInst_MC2_r3Inst_XORInst_0_3_n7,
         MCInst_MC3_v0_2Inst_0_n3, MCInst_MC3_v1_2Inst_0_n3,
         MCInst_MC3_v2_3Inst_0_n6, MCInst_MC3_v2_3Inst_0_n5,
         MCInst_MC3_v3_3Inst_0_n3, MCInst_MC3_v0_2Inst_1_n3,
         MCInst_MC3_v2_1Inst_1_n3, MCInst_MC3_v2_2Inst_1_n6,
         MCInst_MC3_v2_2Inst_1_n5, MCInst_MC3_v3_3Inst_1_n3,
         MCInst_MC3_v1_1Inst_2_n3, MCInst_MC3_v1_2Inst_2_n3,
         MCInst_MC3_v2_1Inst_2_n3, MCInst_MC3_v2_2Inst_2_n3,
         MCInst_MC3_v3_1Inst_2_n3, MCInst_MC3_v1_2Inst_3_n6,
         MCInst_MC3_v1_2Inst_3_n5, MCInst_MC3_v2_2Inst_3_n3,
         MCInst_MC3_v2_3Inst_3_n3, MCInst_MC3_r0Inst_XORInst_0_0_n8,
         MCInst_MC3_r0Inst_XORInst_0_0_n7, MCInst_MC3_r0Inst_XORInst_0_1_n8,
         MCInst_MC3_r0Inst_XORInst_0_1_n7, MCInst_MC3_r0Inst_XORInst_0_2_n8,
         MCInst_MC3_r0Inst_XORInst_0_2_n7, MCInst_MC3_r0Inst_XORInst_0_3_n8,
         MCInst_MC3_r0Inst_XORInst_0_3_n7, MCInst_MC3_r1Inst_XORInst_0_0_n8,
         MCInst_MC3_r1Inst_XORInst_0_0_n7, MCInst_MC3_r1Inst_XORInst_0_1_n8,
         MCInst_MC3_r1Inst_XORInst_0_1_n7, MCInst_MC3_r1Inst_XORInst_0_2_n8,
         MCInst_MC3_r1Inst_XORInst_0_2_n7, MCInst_MC3_r1Inst_XORInst_0_3_n8,
         MCInst_MC3_r1Inst_XORInst_0_3_n7, MCInst_MC3_r2Inst_XORInst_0_0_n8,
         MCInst_MC3_r2Inst_XORInst_0_0_n7, MCInst_MC3_r2Inst_XORInst_0_1_n8,
         MCInst_MC3_r2Inst_XORInst_0_1_n7, MCInst_MC3_r2Inst_XORInst_0_2_n8,
         MCInst_MC3_r2Inst_XORInst_0_2_n7, MCInst_MC3_r2Inst_XORInst_0_3_n8,
         MCInst_MC3_r2Inst_XORInst_0_3_n7, MCInst_MC3_r3Inst_XORInst_0_0_n8,
         MCInst_MC3_r3Inst_XORInst_0_0_n7, MCInst_MC3_r3Inst_XORInst_0_1_n8,
         MCInst_MC3_r3Inst_XORInst_0_1_n7, MCInst_MC3_r3Inst_XORInst_0_2_n8,
         MCInst_MC3_r3Inst_XORInst_0_2_n7, MCInst_MC3_r3Inst_XORInst_0_3_n8,
         MCInst_MC3_r3Inst_XORInst_0_3_n7, SubCellInst2_LFInst_0_LFInst_0_n7,
         SubCellInst2_LFInst_0_LFInst_0_n6, SubCellInst2_LFInst_0_LFInst_0_n5,
         SubCellInst2_LFInst_0_LFInst_1_n26,
         SubCellInst2_LFInst_0_LFInst_1_n25,
         SubCellInst2_LFInst_0_LFInst_1_n24,
         SubCellInst2_LFInst_0_LFInst_1_n23,
         SubCellInst2_LFInst_0_LFInst_1_n22,
         SubCellInst2_LFInst_0_LFInst_1_n21,
         SubCellInst2_LFInst_0_LFInst_1_n20,
         SubCellInst2_LFInst_0_LFInst_1_n19,
         SubCellInst2_LFInst_0_LFInst_1_n18,
         SubCellInst2_LFInst_0_LFInst_2_n28,
         SubCellInst2_LFInst_0_LFInst_2_n27,
         SubCellInst2_LFInst_0_LFInst_2_n26,
         SubCellInst2_LFInst_0_LFInst_2_n25,
         SubCellInst2_LFInst_0_LFInst_2_n24,
         SubCellInst2_LFInst_0_LFInst_2_n23,
         SubCellInst2_LFInst_0_LFInst_2_n22,
         SubCellInst2_LFInst_0_LFInst_3_n26,
         SubCellInst2_LFInst_0_LFInst_3_n25,
         SubCellInst2_LFInst_0_LFInst_3_n24,
         SubCellInst2_LFInst_0_LFInst_3_n23,
         SubCellInst2_LFInst_0_LFInst_3_n22,
         SubCellInst2_LFInst_0_LFInst_3_n21,
         SubCellInst2_LFInst_0_LFInst_3_n20,
         SubCellInst2_LFInst_0_LFInst_3_n19, SubCellInst2_LFInst_1_LFInst_0_n7,
         SubCellInst2_LFInst_1_LFInst_0_n6, SubCellInst2_LFInst_1_LFInst_0_n5,
         SubCellInst2_LFInst_1_LFInst_1_n26,
         SubCellInst2_LFInst_1_LFInst_1_n25,
         SubCellInst2_LFInst_1_LFInst_1_n24,
         SubCellInst2_LFInst_1_LFInst_1_n23,
         SubCellInst2_LFInst_1_LFInst_1_n22,
         SubCellInst2_LFInst_1_LFInst_1_n21,
         SubCellInst2_LFInst_1_LFInst_1_n20,
         SubCellInst2_LFInst_1_LFInst_1_n19,
         SubCellInst2_LFInst_1_LFInst_1_n18,
         SubCellInst2_LFInst_1_LFInst_2_n28,
         SubCellInst2_LFInst_1_LFInst_2_n27,
         SubCellInst2_LFInst_1_LFInst_2_n26,
         SubCellInst2_LFInst_1_LFInst_2_n25,
         SubCellInst2_LFInst_1_LFInst_2_n24,
         SubCellInst2_LFInst_1_LFInst_2_n23,
         SubCellInst2_LFInst_1_LFInst_2_n22,
         SubCellInst2_LFInst_1_LFInst_3_n26,
         SubCellInst2_LFInst_1_LFInst_3_n25,
         SubCellInst2_LFInst_1_LFInst_3_n24,
         SubCellInst2_LFInst_1_LFInst_3_n23,
         SubCellInst2_LFInst_1_LFInst_3_n22,
         SubCellInst2_LFInst_1_LFInst_3_n21,
         SubCellInst2_LFInst_1_LFInst_3_n20,
         SubCellInst2_LFInst_1_LFInst_3_n19, SubCellInst2_LFInst_2_LFInst_0_n7,
         SubCellInst2_LFInst_2_LFInst_0_n6, SubCellInst2_LFInst_2_LFInst_0_n5,
         SubCellInst2_LFInst_2_LFInst_1_n26,
         SubCellInst2_LFInst_2_LFInst_1_n25,
         SubCellInst2_LFInst_2_LFInst_1_n24,
         SubCellInst2_LFInst_2_LFInst_1_n23,
         SubCellInst2_LFInst_2_LFInst_1_n22,
         SubCellInst2_LFInst_2_LFInst_1_n21,
         SubCellInst2_LFInst_2_LFInst_1_n20,
         SubCellInst2_LFInst_2_LFInst_1_n19,
         SubCellInst2_LFInst_2_LFInst_1_n18,
         SubCellInst2_LFInst_2_LFInst_2_n28,
         SubCellInst2_LFInst_2_LFInst_2_n27,
         SubCellInst2_LFInst_2_LFInst_2_n26,
         SubCellInst2_LFInst_2_LFInst_2_n25,
         SubCellInst2_LFInst_2_LFInst_2_n24,
         SubCellInst2_LFInst_2_LFInst_2_n23,
         SubCellInst2_LFInst_2_LFInst_2_n22,
         SubCellInst2_LFInst_2_LFInst_3_n26,
         SubCellInst2_LFInst_2_LFInst_3_n25,
         SubCellInst2_LFInst_2_LFInst_3_n24,
         SubCellInst2_LFInst_2_LFInst_3_n23,
         SubCellInst2_LFInst_2_LFInst_3_n22,
         SubCellInst2_LFInst_2_LFInst_3_n21,
         SubCellInst2_LFInst_2_LFInst_3_n20,
         SubCellInst2_LFInst_2_LFInst_3_n19, SubCellInst2_LFInst_3_LFInst_0_n7,
         SubCellInst2_LFInst_3_LFInst_0_n6, SubCellInst2_LFInst_3_LFInst_0_n5,
         SubCellInst2_LFInst_3_LFInst_1_n26,
         SubCellInst2_LFInst_3_LFInst_1_n25,
         SubCellInst2_LFInst_3_LFInst_1_n24,
         SubCellInst2_LFInst_3_LFInst_1_n23,
         SubCellInst2_LFInst_3_LFInst_1_n22,
         SubCellInst2_LFInst_3_LFInst_1_n21,
         SubCellInst2_LFInst_3_LFInst_1_n20,
         SubCellInst2_LFInst_3_LFInst_1_n19,
         SubCellInst2_LFInst_3_LFInst_1_n18,
         SubCellInst2_LFInst_3_LFInst_2_n28,
         SubCellInst2_LFInst_3_LFInst_2_n27,
         SubCellInst2_LFInst_3_LFInst_2_n26,
         SubCellInst2_LFInst_3_LFInst_2_n25,
         SubCellInst2_LFInst_3_LFInst_2_n24,
         SubCellInst2_LFInst_3_LFInst_2_n23,
         SubCellInst2_LFInst_3_LFInst_2_n22,
         SubCellInst2_LFInst_3_LFInst_3_n26,
         SubCellInst2_LFInst_3_LFInst_3_n25,
         SubCellInst2_LFInst_3_LFInst_3_n24,
         SubCellInst2_LFInst_3_LFInst_3_n23,
         SubCellInst2_LFInst_3_LFInst_3_n22,
         SubCellInst2_LFInst_3_LFInst_3_n21,
         SubCellInst2_LFInst_3_LFInst_3_n20,
         SubCellInst2_LFInst_3_LFInst_3_n19, SubCellInst2_LFInst_4_LFInst_0_n7,
         SubCellInst2_LFInst_4_LFInst_0_n6, SubCellInst2_LFInst_4_LFInst_0_n5,
         SubCellInst2_LFInst_4_LFInst_1_n26,
         SubCellInst2_LFInst_4_LFInst_1_n25,
         SubCellInst2_LFInst_4_LFInst_1_n24,
         SubCellInst2_LFInst_4_LFInst_1_n23,
         SubCellInst2_LFInst_4_LFInst_1_n22,
         SubCellInst2_LFInst_4_LFInst_1_n21,
         SubCellInst2_LFInst_4_LFInst_1_n20,
         SubCellInst2_LFInst_4_LFInst_1_n19,
         SubCellInst2_LFInst_4_LFInst_1_n18,
         SubCellInst2_LFInst_4_LFInst_2_n29,
         SubCellInst2_LFInst_4_LFInst_2_n28,
         SubCellInst2_LFInst_4_LFInst_2_n27,
         SubCellInst2_LFInst_4_LFInst_2_n26,
         SubCellInst2_LFInst_4_LFInst_2_n25,
         SubCellInst2_LFInst_4_LFInst_2_n24,
         SubCellInst2_LFInst_4_LFInst_2_n23,
         SubCellInst2_LFInst_4_LFInst_2_n22,
         SubCellInst2_LFInst_4_LFInst_3_n26,
         SubCellInst2_LFInst_4_LFInst_3_n25,
         SubCellInst2_LFInst_4_LFInst_3_n24,
         SubCellInst2_LFInst_4_LFInst_3_n23,
         SubCellInst2_LFInst_4_LFInst_3_n22,
         SubCellInst2_LFInst_4_LFInst_3_n21,
         SubCellInst2_LFInst_4_LFInst_3_n20,
         SubCellInst2_LFInst_4_LFInst_3_n19, SubCellInst2_LFInst_5_LFInst_0_n7,
         SubCellInst2_LFInst_5_LFInst_0_n6, SubCellInst2_LFInst_5_LFInst_0_n5,
         SubCellInst2_LFInst_5_LFInst_1_n26,
         SubCellInst2_LFInst_5_LFInst_1_n25,
         SubCellInst2_LFInst_5_LFInst_1_n24,
         SubCellInst2_LFInst_5_LFInst_1_n23,
         SubCellInst2_LFInst_5_LFInst_1_n22,
         SubCellInst2_LFInst_5_LFInst_1_n21,
         SubCellInst2_LFInst_5_LFInst_1_n20,
         SubCellInst2_LFInst_5_LFInst_1_n19,
         SubCellInst2_LFInst_5_LFInst_1_n18,
         SubCellInst2_LFInst_5_LFInst_2_n29,
         SubCellInst2_LFInst_5_LFInst_2_n28,
         SubCellInst2_LFInst_5_LFInst_2_n27,
         SubCellInst2_LFInst_5_LFInst_2_n26,
         SubCellInst2_LFInst_5_LFInst_2_n25,
         SubCellInst2_LFInst_5_LFInst_2_n24,
         SubCellInst2_LFInst_5_LFInst_2_n23,
         SubCellInst2_LFInst_5_LFInst_2_n22,
         SubCellInst2_LFInst_5_LFInst_3_n26,
         SubCellInst2_LFInst_5_LFInst_3_n25,
         SubCellInst2_LFInst_5_LFInst_3_n24,
         SubCellInst2_LFInst_5_LFInst_3_n23,
         SubCellInst2_LFInst_5_LFInst_3_n22,
         SubCellInst2_LFInst_5_LFInst_3_n21,
         SubCellInst2_LFInst_5_LFInst_3_n20,
         SubCellInst2_LFInst_5_LFInst_3_n19, SubCellInst2_LFInst_6_LFInst_0_n7,
         SubCellInst2_LFInst_6_LFInst_0_n6, SubCellInst2_LFInst_6_LFInst_0_n5,
         SubCellInst2_LFInst_6_LFInst_1_n26,
         SubCellInst2_LFInst_6_LFInst_1_n25,
         SubCellInst2_LFInst_6_LFInst_1_n24,
         SubCellInst2_LFInst_6_LFInst_1_n23,
         SubCellInst2_LFInst_6_LFInst_1_n22,
         SubCellInst2_LFInst_6_LFInst_1_n21,
         SubCellInst2_LFInst_6_LFInst_1_n20,
         SubCellInst2_LFInst_6_LFInst_1_n19,
         SubCellInst2_LFInst_6_LFInst_1_n18,
         SubCellInst2_LFInst_6_LFInst_2_n29,
         SubCellInst2_LFInst_6_LFInst_2_n28,
         SubCellInst2_LFInst_6_LFInst_2_n27,
         SubCellInst2_LFInst_6_LFInst_2_n26,
         SubCellInst2_LFInst_6_LFInst_2_n25,
         SubCellInst2_LFInst_6_LFInst_2_n24,
         SubCellInst2_LFInst_6_LFInst_2_n23,
         SubCellInst2_LFInst_6_LFInst_2_n22,
         SubCellInst2_LFInst_6_LFInst_3_n26,
         SubCellInst2_LFInst_6_LFInst_3_n25,
         SubCellInst2_LFInst_6_LFInst_3_n24,
         SubCellInst2_LFInst_6_LFInst_3_n23,
         SubCellInst2_LFInst_6_LFInst_3_n22,
         SubCellInst2_LFInst_6_LFInst_3_n21,
         SubCellInst2_LFInst_6_LFInst_3_n20,
         SubCellInst2_LFInst_6_LFInst_3_n19, SubCellInst2_LFInst_7_LFInst_0_n7,
         SubCellInst2_LFInst_7_LFInst_0_n6, SubCellInst2_LFInst_7_LFInst_0_n5,
         SubCellInst2_LFInst_7_LFInst_1_n26,
         SubCellInst2_LFInst_7_LFInst_1_n25,
         SubCellInst2_LFInst_7_LFInst_1_n24,
         SubCellInst2_LFInst_7_LFInst_1_n23,
         SubCellInst2_LFInst_7_LFInst_1_n22,
         SubCellInst2_LFInst_7_LFInst_1_n21,
         SubCellInst2_LFInst_7_LFInst_1_n20,
         SubCellInst2_LFInst_7_LFInst_1_n19,
         SubCellInst2_LFInst_7_LFInst_1_n18,
         SubCellInst2_LFInst_7_LFInst_2_n29,
         SubCellInst2_LFInst_7_LFInst_2_n28,
         SubCellInst2_LFInst_7_LFInst_2_n27,
         SubCellInst2_LFInst_7_LFInst_2_n26,
         SubCellInst2_LFInst_7_LFInst_2_n25,
         SubCellInst2_LFInst_7_LFInst_2_n24,
         SubCellInst2_LFInst_7_LFInst_2_n23,
         SubCellInst2_LFInst_7_LFInst_2_n22,
         SubCellInst2_LFInst_7_LFInst_3_n26,
         SubCellInst2_LFInst_7_LFInst_3_n25,
         SubCellInst2_LFInst_7_LFInst_3_n24,
         SubCellInst2_LFInst_7_LFInst_3_n23,
         SubCellInst2_LFInst_7_LFInst_3_n22,
         SubCellInst2_LFInst_7_LFInst_3_n21,
         SubCellInst2_LFInst_7_LFInst_3_n20,
         SubCellInst2_LFInst_7_LFInst_3_n19, SubCellInst2_LFInst_8_LFInst_0_n7,
         SubCellInst2_LFInst_8_LFInst_0_n6, SubCellInst2_LFInst_8_LFInst_0_n5,
         SubCellInst2_LFInst_8_LFInst_1_n26,
         SubCellInst2_LFInst_8_LFInst_1_n25,
         SubCellInst2_LFInst_8_LFInst_1_n24,
         SubCellInst2_LFInst_8_LFInst_1_n23,
         SubCellInst2_LFInst_8_LFInst_1_n22,
         SubCellInst2_LFInst_8_LFInst_1_n21,
         SubCellInst2_LFInst_8_LFInst_1_n20,
         SubCellInst2_LFInst_8_LFInst_1_n19,
         SubCellInst2_LFInst_8_LFInst_1_n18,
         SubCellInst2_LFInst_8_LFInst_2_n29,
         SubCellInst2_LFInst_8_LFInst_2_n28,
         SubCellInst2_LFInst_8_LFInst_2_n27,
         SubCellInst2_LFInst_8_LFInst_2_n26,
         SubCellInst2_LFInst_8_LFInst_2_n25,
         SubCellInst2_LFInst_8_LFInst_2_n24,
         SubCellInst2_LFInst_8_LFInst_2_n23,
         SubCellInst2_LFInst_8_LFInst_2_n22,
         SubCellInst2_LFInst_8_LFInst_3_n26,
         SubCellInst2_LFInst_8_LFInst_3_n25,
         SubCellInst2_LFInst_8_LFInst_3_n24,
         SubCellInst2_LFInst_8_LFInst_3_n23,
         SubCellInst2_LFInst_8_LFInst_3_n22,
         SubCellInst2_LFInst_8_LFInst_3_n21,
         SubCellInst2_LFInst_8_LFInst_3_n20,
         SubCellInst2_LFInst_8_LFInst_3_n19, SubCellInst2_LFInst_9_LFInst_0_n7,
         SubCellInst2_LFInst_9_LFInst_0_n6, SubCellInst2_LFInst_9_LFInst_0_n5,
         SubCellInst2_LFInst_9_LFInst_1_n26,
         SubCellInst2_LFInst_9_LFInst_1_n25,
         SubCellInst2_LFInst_9_LFInst_1_n24,
         SubCellInst2_LFInst_9_LFInst_1_n23,
         SubCellInst2_LFInst_9_LFInst_1_n22,
         SubCellInst2_LFInst_9_LFInst_1_n21,
         SubCellInst2_LFInst_9_LFInst_1_n20,
         SubCellInst2_LFInst_9_LFInst_1_n19,
         SubCellInst2_LFInst_9_LFInst_1_n18,
         SubCellInst2_LFInst_9_LFInst_2_n29,
         SubCellInst2_LFInst_9_LFInst_2_n28,
         SubCellInst2_LFInst_9_LFInst_2_n27,
         SubCellInst2_LFInst_9_LFInst_2_n26,
         SubCellInst2_LFInst_9_LFInst_2_n25,
         SubCellInst2_LFInst_9_LFInst_2_n24,
         SubCellInst2_LFInst_9_LFInst_2_n23,
         SubCellInst2_LFInst_9_LFInst_2_n22,
         SubCellInst2_LFInst_9_LFInst_3_n26,
         SubCellInst2_LFInst_9_LFInst_3_n25,
         SubCellInst2_LFInst_9_LFInst_3_n24,
         SubCellInst2_LFInst_9_LFInst_3_n23,
         SubCellInst2_LFInst_9_LFInst_3_n22,
         SubCellInst2_LFInst_9_LFInst_3_n21,
         SubCellInst2_LFInst_9_LFInst_3_n20,
         SubCellInst2_LFInst_9_LFInst_3_n19,
         SubCellInst2_LFInst_10_LFInst_0_n7,
         SubCellInst2_LFInst_10_LFInst_0_n6,
         SubCellInst2_LFInst_10_LFInst_0_n5,
         SubCellInst2_LFInst_10_LFInst_1_n26,
         SubCellInst2_LFInst_10_LFInst_1_n25,
         SubCellInst2_LFInst_10_LFInst_1_n24,
         SubCellInst2_LFInst_10_LFInst_1_n23,
         SubCellInst2_LFInst_10_LFInst_1_n22,
         SubCellInst2_LFInst_10_LFInst_1_n21,
         SubCellInst2_LFInst_10_LFInst_1_n20,
         SubCellInst2_LFInst_10_LFInst_1_n19,
         SubCellInst2_LFInst_10_LFInst_1_n18,
         SubCellInst2_LFInst_10_LFInst_2_n29,
         SubCellInst2_LFInst_10_LFInst_2_n28,
         SubCellInst2_LFInst_10_LFInst_2_n27,
         SubCellInst2_LFInst_10_LFInst_2_n26,
         SubCellInst2_LFInst_10_LFInst_2_n25,
         SubCellInst2_LFInst_10_LFInst_2_n24,
         SubCellInst2_LFInst_10_LFInst_2_n23,
         SubCellInst2_LFInst_10_LFInst_2_n22,
         SubCellInst2_LFInst_10_LFInst_3_n26,
         SubCellInst2_LFInst_10_LFInst_3_n25,
         SubCellInst2_LFInst_10_LFInst_3_n24,
         SubCellInst2_LFInst_10_LFInst_3_n23,
         SubCellInst2_LFInst_10_LFInst_3_n22,
         SubCellInst2_LFInst_10_LFInst_3_n21,
         SubCellInst2_LFInst_10_LFInst_3_n20,
         SubCellInst2_LFInst_10_LFInst_3_n19,
         SubCellInst2_LFInst_11_LFInst_0_n7,
         SubCellInst2_LFInst_11_LFInst_0_n6,
         SubCellInst2_LFInst_11_LFInst_0_n5,
         SubCellInst2_LFInst_11_LFInst_1_n26,
         SubCellInst2_LFInst_11_LFInst_1_n25,
         SubCellInst2_LFInst_11_LFInst_1_n24,
         SubCellInst2_LFInst_11_LFInst_1_n23,
         SubCellInst2_LFInst_11_LFInst_1_n22,
         SubCellInst2_LFInst_11_LFInst_1_n21,
         SubCellInst2_LFInst_11_LFInst_1_n20,
         SubCellInst2_LFInst_11_LFInst_1_n19,
         SubCellInst2_LFInst_11_LFInst_1_n18,
         SubCellInst2_LFInst_11_LFInst_2_n29,
         SubCellInst2_LFInst_11_LFInst_2_n28,
         SubCellInst2_LFInst_11_LFInst_2_n27,
         SubCellInst2_LFInst_11_LFInst_2_n26,
         SubCellInst2_LFInst_11_LFInst_2_n25,
         SubCellInst2_LFInst_11_LFInst_2_n24,
         SubCellInst2_LFInst_11_LFInst_2_n23,
         SubCellInst2_LFInst_11_LFInst_2_n22,
         SubCellInst2_LFInst_11_LFInst_3_n26,
         SubCellInst2_LFInst_11_LFInst_3_n25,
         SubCellInst2_LFInst_11_LFInst_3_n24,
         SubCellInst2_LFInst_11_LFInst_3_n23,
         SubCellInst2_LFInst_11_LFInst_3_n22,
         SubCellInst2_LFInst_11_LFInst_3_n21,
         SubCellInst2_LFInst_11_LFInst_3_n20,
         SubCellInst2_LFInst_11_LFInst_3_n19,
         SubCellInst2_LFInst_12_LFInst_0_n7,
         SubCellInst2_LFInst_12_LFInst_0_n6,
         SubCellInst2_LFInst_12_LFInst_0_n5,
         SubCellInst2_LFInst_12_LFInst_1_n26,
         SubCellInst2_LFInst_12_LFInst_1_n25,
         SubCellInst2_LFInst_12_LFInst_1_n24,
         SubCellInst2_LFInst_12_LFInst_1_n23,
         SubCellInst2_LFInst_12_LFInst_1_n22,
         SubCellInst2_LFInst_12_LFInst_1_n21,
         SubCellInst2_LFInst_12_LFInst_1_n20,
         SubCellInst2_LFInst_12_LFInst_1_n19,
         SubCellInst2_LFInst_12_LFInst_1_n18,
         SubCellInst2_LFInst_12_LFInst_2_n29,
         SubCellInst2_LFInst_12_LFInst_2_n28,
         SubCellInst2_LFInst_12_LFInst_2_n27,
         SubCellInst2_LFInst_12_LFInst_2_n26,
         SubCellInst2_LFInst_12_LFInst_2_n25,
         SubCellInst2_LFInst_12_LFInst_2_n24,
         SubCellInst2_LFInst_12_LFInst_2_n23,
         SubCellInst2_LFInst_12_LFInst_2_n22,
         SubCellInst2_LFInst_12_LFInst_3_n26,
         SubCellInst2_LFInst_12_LFInst_3_n25,
         SubCellInst2_LFInst_12_LFInst_3_n24,
         SubCellInst2_LFInst_12_LFInst_3_n23,
         SubCellInst2_LFInst_12_LFInst_3_n22,
         SubCellInst2_LFInst_12_LFInst_3_n21,
         SubCellInst2_LFInst_12_LFInst_3_n20,
         SubCellInst2_LFInst_12_LFInst_3_n19,
         SubCellInst2_LFInst_13_LFInst_0_n7,
         SubCellInst2_LFInst_13_LFInst_0_n6,
         SubCellInst2_LFInst_13_LFInst_0_n5,
         SubCellInst2_LFInst_13_LFInst_1_n26,
         SubCellInst2_LFInst_13_LFInst_1_n25,
         SubCellInst2_LFInst_13_LFInst_1_n24,
         SubCellInst2_LFInst_13_LFInst_1_n23,
         SubCellInst2_LFInst_13_LFInst_1_n22,
         SubCellInst2_LFInst_13_LFInst_1_n21,
         SubCellInst2_LFInst_13_LFInst_1_n20,
         SubCellInst2_LFInst_13_LFInst_1_n19,
         SubCellInst2_LFInst_13_LFInst_1_n18,
         SubCellInst2_LFInst_13_LFInst_2_n29,
         SubCellInst2_LFInst_13_LFInst_2_n28,
         SubCellInst2_LFInst_13_LFInst_2_n27,
         SubCellInst2_LFInst_13_LFInst_2_n26,
         SubCellInst2_LFInst_13_LFInst_2_n25,
         SubCellInst2_LFInst_13_LFInst_2_n24,
         SubCellInst2_LFInst_13_LFInst_2_n23,
         SubCellInst2_LFInst_13_LFInst_2_n22,
         SubCellInst2_LFInst_13_LFInst_3_n26,
         SubCellInst2_LFInst_13_LFInst_3_n25,
         SubCellInst2_LFInst_13_LFInst_3_n24,
         SubCellInst2_LFInst_13_LFInst_3_n23,
         SubCellInst2_LFInst_13_LFInst_3_n22,
         SubCellInst2_LFInst_13_LFInst_3_n21,
         SubCellInst2_LFInst_13_LFInst_3_n20,
         SubCellInst2_LFInst_13_LFInst_3_n19,
         SubCellInst2_LFInst_14_LFInst_0_n7,
         SubCellInst2_LFInst_14_LFInst_0_n6,
         SubCellInst2_LFInst_14_LFInst_0_n5,
         SubCellInst2_LFInst_14_LFInst_1_n26,
         SubCellInst2_LFInst_14_LFInst_1_n25,
         SubCellInst2_LFInst_14_LFInst_1_n24,
         SubCellInst2_LFInst_14_LFInst_1_n23,
         SubCellInst2_LFInst_14_LFInst_1_n22,
         SubCellInst2_LFInst_14_LFInst_1_n21,
         SubCellInst2_LFInst_14_LFInst_1_n20,
         SubCellInst2_LFInst_14_LFInst_1_n19,
         SubCellInst2_LFInst_14_LFInst_1_n18,
         SubCellInst2_LFInst_14_LFInst_2_n29,
         SubCellInst2_LFInst_14_LFInst_2_n28,
         SubCellInst2_LFInst_14_LFInst_2_n27,
         SubCellInst2_LFInst_14_LFInst_2_n26,
         SubCellInst2_LFInst_14_LFInst_2_n25,
         SubCellInst2_LFInst_14_LFInst_2_n24,
         SubCellInst2_LFInst_14_LFInst_2_n23,
         SubCellInst2_LFInst_14_LFInst_2_n22,
         SubCellInst2_LFInst_14_LFInst_3_n26,
         SubCellInst2_LFInst_14_LFInst_3_n25,
         SubCellInst2_LFInst_14_LFInst_3_n24,
         SubCellInst2_LFInst_14_LFInst_3_n23,
         SubCellInst2_LFInst_14_LFInst_3_n22,
         SubCellInst2_LFInst_14_LFInst_3_n21,
         SubCellInst2_LFInst_14_LFInst_3_n20,
         SubCellInst2_LFInst_14_LFInst_3_n19,
         SubCellInst2_LFInst_15_LFInst_0_n7,
         SubCellInst2_LFInst_15_LFInst_0_n6,
         SubCellInst2_LFInst_15_LFInst_0_n5,
         SubCellInst2_LFInst_15_LFInst_1_n26,
         SubCellInst2_LFInst_15_LFInst_1_n25,
         SubCellInst2_LFInst_15_LFInst_1_n24,
         SubCellInst2_LFInst_15_LFInst_1_n23,
         SubCellInst2_LFInst_15_LFInst_1_n22,
         SubCellInst2_LFInst_15_LFInst_1_n21,
         SubCellInst2_LFInst_15_LFInst_1_n20,
         SubCellInst2_LFInst_15_LFInst_1_n19,
         SubCellInst2_LFInst_15_LFInst_1_n18,
         SubCellInst2_LFInst_15_LFInst_2_n29,
         SubCellInst2_LFInst_15_LFInst_2_n28,
         SubCellInst2_LFInst_15_LFInst_2_n27,
         SubCellInst2_LFInst_15_LFInst_2_n26,
         SubCellInst2_LFInst_15_LFInst_2_n25,
         SubCellInst2_LFInst_15_LFInst_2_n24,
         SubCellInst2_LFInst_15_LFInst_2_n23,
         SubCellInst2_LFInst_15_LFInst_2_n22,
         SubCellInst2_LFInst_15_LFInst_3_n26,
         SubCellInst2_LFInst_15_LFInst_3_n25,
         SubCellInst2_LFInst_15_LFInst_3_n24,
         SubCellInst2_LFInst_15_LFInst_3_n23,
         SubCellInst2_LFInst_15_LFInst_3_n22,
         SubCellInst2_LFInst_15_LFInst_3_n21,
         SubCellInst2_LFInst_15_LFInst_3_n20,
         SubCellInst2_LFInst_15_LFInst_3_n19, MCInst2_MC0_v0_2Inst_0_n3,
         MCInst2_MC0_v1_2Inst_0_n3, MCInst2_MC0_v2_3Inst_0_n6,
         MCInst2_MC0_v2_3Inst_0_n5, MCInst2_MC0_v3_3Inst_0_n3,
         MCInst2_MC0_v0_2Inst_1_n3, MCInst2_MC0_v2_1Inst_1_n3,
         MCInst2_MC0_v2_2Inst_1_n6, MCInst2_MC0_v2_2Inst_1_n5,
         MCInst2_MC0_v3_3Inst_1_n3, MCInst2_MC0_v1_1Inst_2_n3,
         MCInst2_MC0_v1_2Inst_2_n3, MCInst2_MC0_v2_1Inst_2_n3,
         MCInst2_MC0_v2_2Inst_2_n3, MCInst2_MC0_v3_1Inst_2_n3,
         MCInst2_MC0_v1_2Inst_3_n6, MCInst2_MC0_v1_2Inst_3_n5,
         MCInst2_MC0_v2_2Inst_3_n3, MCInst2_MC0_v2_3Inst_3_n3,
         MCInst2_MC0_r0Inst_XORInst_0_0_n8, MCInst2_MC0_r0Inst_XORInst_0_0_n7,
         MCInst2_MC0_r0Inst_XORInst_0_1_n8, MCInst2_MC0_r0Inst_XORInst_0_1_n7,
         MCInst2_MC0_r0Inst_XORInst_0_2_n8, MCInst2_MC0_r0Inst_XORInst_0_2_n7,
         MCInst2_MC0_r0Inst_XORInst_0_3_n8, MCInst2_MC0_r0Inst_XORInst_0_3_n7,
         MCInst2_MC0_r1Inst_XORInst_0_0_n8, MCInst2_MC0_r1Inst_XORInst_0_0_n7,
         MCInst2_MC0_r1Inst_XORInst_0_1_n8, MCInst2_MC0_r1Inst_XORInst_0_1_n7,
         MCInst2_MC0_r1Inst_XORInst_0_2_n8, MCInst2_MC0_r1Inst_XORInst_0_2_n7,
         MCInst2_MC0_r1Inst_XORInst_0_3_n8, MCInst2_MC0_r1Inst_XORInst_0_3_n7,
         MCInst2_MC0_r2Inst_XORInst_0_0_n8, MCInst2_MC0_r2Inst_XORInst_0_0_n7,
         MCInst2_MC0_r2Inst_XORInst_0_1_n8, MCInst2_MC0_r2Inst_XORInst_0_1_n7,
         MCInst2_MC0_r2Inst_XORInst_0_2_n8, MCInst2_MC0_r2Inst_XORInst_0_2_n7,
         MCInst2_MC0_r2Inst_XORInst_0_3_n8, MCInst2_MC0_r2Inst_XORInst_0_3_n7,
         MCInst2_MC0_r3Inst_XORInst_0_0_n8, MCInst2_MC0_r3Inst_XORInst_0_0_n7,
         MCInst2_MC0_r3Inst_XORInst_0_1_n8, MCInst2_MC0_r3Inst_XORInst_0_1_n7,
         MCInst2_MC0_r3Inst_XORInst_0_2_n8, MCInst2_MC0_r3Inst_XORInst_0_2_n7,
         MCInst2_MC0_r3Inst_XORInst_0_3_n8, MCInst2_MC0_r3Inst_XORInst_0_3_n7,
         MCInst2_MC1_v0_2Inst_0_n3, MCInst2_MC1_v1_2Inst_0_n3,
         MCInst2_MC1_v2_3Inst_0_n6, MCInst2_MC1_v2_3Inst_0_n5,
         MCInst2_MC1_v3_3Inst_0_n3, MCInst2_MC1_v0_2Inst_1_n3,
         MCInst2_MC1_v2_1Inst_1_n3, MCInst2_MC1_v2_2Inst_1_n6,
         MCInst2_MC1_v2_2Inst_1_n5, MCInst2_MC1_v3_3Inst_1_n3,
         MCInst2_MC1_v1_1Inst_2_n3, MCInst2_MC1_v1_2Inst_2_n3,
         MCInst2_MC1_v2_1Inst_2_n3, MCInst2_MC1_v2_2Inst_2_n3,
         MCInst2_MC1_v3_1Inst_2_n3, MCInst2_MC1_v1_2Inst_3_n6,
         MCInst2_MC1_v1_2Inst_3_n5, MCInst2_MC1_v2_2Inst_3_n3,
         MCInst2_MC1_v2_3Inst_3_n3, MCInst2_MC1_r0Inst_XORInst_0_0_n8,
         MCInst2_MC1_r0Inst_XORInst_0_0_n7, MCInst2_MC1_r0Inst_XORInst_0_1_n8,
         MCInst2_MC1_r0Inst_XORInst_0_1_n7, MCInst2_MC1_r0Inst_XORInst_0_2_n8,
         MCInst2_MC1_r0Inst_XORInst_0_2_n7, MCInst2_MC1_r0Inst_XORInst_0_3_n8,
         MCInst2_MC1_r0Inst_XORInst_0_3_n7, MCInst2_MC1_r1Inst_XORInst_0_0_n8,
         MCInst2_MC1_r1Inst_XORInst_0_0_n7, MCInst2_MC1_r1Inst_XORInst_0_1_n8,
         MCInst2_MC1_r1Inst_XORInst_0_1_n7, MCInst2_MC1_r1Inst_XORInst_0_2_n8,
         MCInst2_MC1_r1Inst_XORInst_0_2_n7, MCInst2_MC1_r1Inst_XORInst_0_3_n8,
         MCInst2_MC1_r1Inst_XORInst_0_3_n7, MCInst2_MC1_r2Inst_XORInst_0_0_n8,
         MCInst2_MC1_r2Inst_XORInst_0_0_n7, MCInst2_MC1_r2Inst_XORInst_0_1_n8,
         MCInst2_MC1_r2Inst_XORInst_0_1_n7, MCInst2_MC1_r2Inst_XORInst_0_2_n8,
         MCInst2_MC1_r2Inst_XORInst_0_2_n7, MCInst2_MC1_r2Inst_XORInst_0_3_n8,
         MCInst2_MC1_r2Inst_XORInst_0_3_n7, MCInst2_MC1_r3Inst_XORInst_0_0_n8,
         MCInst2_MC1_r3Inst_XORInst_0_0_n7, MCInst2_MC1_r3Inst_XORInst_0_1_n8,
         MCInst2_MC1_r3Inst_XORInst_0_1_n7, MCInst2_MC1_r3Inst_XORInst_0_2_n8,
         MCInst2_MC1_r3Inst_XORInst_0_2_n7, MCInst2_MC1_r3Inst_XORInst_0_3_n8,
         MCInst2_MC1_r3Inst_XORInst_0_3_n7, MCInst2_MC2_v0_2Inst_0_n3,
         MCInst2_MC2_v1_2Inst_0_n3, MCInst2_MC2_v2_3Inst_0_n6,
         MCInst2_MC2_v2_3Inst_0_n5, MCInst2_MC2_v3_3Inst_0_n3,
         MCInst2_MC2_v0_2Inst_1_n3, MCInst2_MC2_v2_1Inst_1_n3,
         MCInst2_MC2_v2_2Inst_1_n6, MCInst2_MC2_v2_2Inst_1_n5,
         MCInst2_MC2_v3_3Inst_1_n3, MCInst2_MC2_v1_1Inst_2_n3,
         MCInst2_MC2_v1_2Inst_2_n3, MCInst2_MC2_v2_1Inst_2_n3,
         MCInst2_MC2_v2_2Inst_2_n3, MCInst2_MC2_v3_1Inst_2_n3,
         MCInst2_MC2_v1_2Inst_3_n6, MCInst2_MC2_v1_2Inst_3_n5,
         MCInst2_MC2_v2_2Inst_3_n3, MCInst2_MC2_v2_3Inst_3_n3,
         MCInst2_MC2_r0Inst_XORInst_0_0_n8, MCInst2_MC2_r0Inst_XORInst_0_0_n7,
         MCInst2_MC2_r0Inst_XORInst_0_1_n8, MCInst2_MC2_r0Inst_XORInst_0_1_n7,
         MCInst2_MC2_r0Inst_XORInst_0_2_n8, MCInst2_MC2_r0Inst_XORInst_0_2_n7,
         MCInst2_MC2_r0Inst_XORInst_0_3_n8, MCInst2_MC2_r0Inst_XORInst_0_3_n7,
         MCInst2_MC2_r1Inst_XORInst_0_0_n8, MCInst2_MC2_r1Inst_XORInst_0_0_n7,
         MCInst2_MC2_r1Inst_XORInst_0_1_n8, MCInst2_MC2_r1Inst_XORInst_0_1_n7,
         MCInst2_MC2_r1Inst_XORInst_0_2_n8, MCInst2_MC2_r1Inst_XORInst_0_2_n7,
         MCInst2_MC2_r1Inst_XORInst_0_3_n8, MCInst2_MC2_r1Inst_XORInst_0_3_n7,
         MCInst2_MC2_r2Inst_XORInst_0_0_n8, MCInst2_MC2_r2Inst_XORInst_0_0_n7,
         MCInst2_MC2_r2Inst_XORInst_0_1_n8, MCInst2_MC2_r2Inst_XORInst_0_1_n7,
         MCInst2_MC2_r2Inst_XORInst_0_2_n8, MCInst2_MC2_r2Inst_XORInst_0_2_n7,
         MCInst2_MC2_r2Inst_XORInst_0_3_n8, MCInst2_MC2_r2Inst_XORInst_0_3_n7,
         MCInst2_MC2_r3Inst_XORInst_0_0_n8, MCInst2_MC2_r3Inst_XORInst_0_0_n7,
         MCInst2_MC2_r3Inst_XORInst_0_1_n8, MCInst2_MC2_r3Inst_XORInst_0_1_n7,
         MCInst2_MC2_r3Inst_XORInst_0_2_n8, MCInst2_MC2_r3Inst_XORInst_0_2_n7,
         MCInst2_MC2_r3Inst_XORInst_0_3_n8, MCInst2_MC2_r3Inst_XORInst_0_3_n7,
         MCInst2_MC3_v0_2Inst_0_n3, MCInst2_MC3_v1_2Inst_0_n3,
         MCInst2_MC3_v2_3Inst_0_n6, MCInst2_MC3_v2_3Inst_0_n5,
         MCInst2_MC3_v3_3Inst_0_n3, MCInst2_MC3_v0_2Inst_1_n3,
         MCInst2_MC3_v2_1Inst_1_n3, MCInst2_MC3_v2_2Inst_1_n6,
         MCInst2_MC3_v2_2Inst_1_n5, MCInst2_MC3_v3_3Inst_1_n3,
         MCInst2_MC3_v1_1Inst_2_n3, MCInst2_MC3_v1_2Inst_2_n3,
         MCInst2_MC3_v2_1Inst_2_n3, MCInst2_MC3_v2_2Inst_2_n3,
         MCInst2_MC3_v3_1Inst_2_n3, MCInst2_MC3_v1_2Inst_3_n6,
         MCInst2_MC3_v1_2Inst_3_n5, MCInst2_MC3_v2_2Inst_3_n3,
         MCInst2_MC3_v2_3Inst_3_n3, MCInst2_MC3_r0Inst_XORInst_0_0_n8,
         MCInst2_MC3_r0Inst_XORInst_0_0_n7, MCInst2_MC3_r0Inst_XORInst_0_1_n8,
         MCInst2_MC3_r0Inst_XORInst_0_1_n7, MCInst2_MC3_r0Inst_XORInst_0_2_n8,
         MCInst2_MC3_r0Inst_XORInst_0_2_n7, MCInst2_MC3_r0Inst_XORInst_0_3_n8,
         MCInst2_MC3_r0Inst_XORInst_0_3_n7, MCInst2_MC3_r1Inst_XORInst_0_0_n8,
         MCInst2_MC3_r1Inst_XORInst_0_0_n7, MCInst2_MC3_r1Inst_XORInst_0_1_n8,
         MCInst2_MC3_r1Inst_XORInst_0_1_n7, MCInst2_MC3_r1Inst_XORInst_0_2_n8,
         MCInst2_MC3_r1Inst_XORInst_0_2_n7, MCInst2_MC3_r1Inst_XORInst_0_3_n8,
         MCInst2_MC3_r1Inst_XORInst_0_3_n7, MCInst2_MC3_r2Inst_XORInst_0_0_n8,
         MCInst2_MC3_r2Inst_XORInst_0_0_n7, MCInst2_MC3_r2Inst_XORInst_0_1_n8,
         MCInst2_MC3_r2Inst_XORInst_0_1_n7, MCInst2_MC3_r2Inst_XORInst_0_2_n8,
         MCInst2_MC3_r2Inst_XORInst_0_2_n7, MCInst2_MC3_r2Inst_XORInst_0_3_n8,
         MCInst2_MC3_r2Inst_XORInst_0_3_n7, MCInst2_MC3_r3Inst_XORInst_0_0_n8,
         MCInst2_MC3_r3Inst_XORInst_0_0_n7, MCInst2_MC3_r3Inst_XORInst_0_1_n8,
         MCInst2_MC3_r3Inst_XORInst_0_1_n7, MCInst2_MC3_r3Inst_XORInst_0_2_n8,
         MCInst2_MC3_r3Inst_XORInst_0_2_n7, MCInst2_MC3_r3Inst_XORInst_0_3_n8,
         MCInst2_MC3_r3Inst_XORInst_0_3_n7,
         Red_PlaintextInst_LFInst_0_LFInst_0_n6,
         Red_PlaintextInst_LFInst_0_LFInst_0_n5,
         Red_PlaintextInst_LFInst_1_LFInst_0_n6,
         Red_PlaintextInst_LFInst_1_LFInst_0_n5,
         Red_PlaintextInst_LFInst_2_LFInst_0_n6,
         Red_PlaintextInst_LFInst_2_LFInst_0_n5,
         Red_PlaintextInst_LFInst_3_LFInst_0_n6,
         Red_PlaintextInst_LFInst_3_LFInst_0_n5,
         Red_PlaintextInst_LFInst_4_LFInst_0_n6,
         Red_PlaintextInst_LFInst_4_LFInst_0_n5,
         Red_PlaintextInst_LFInst_5_LFInst_0_n6,
         Red_PlaintextInst_LFInst_5_LFInst_0_n5,
         Red_PlaintextInst_LFInst_6_LFInst_0_n6,
         Red_PlaintextInst_LFInst_6_LFInst_0_n5,
         Red_PlaintextInst_LFInst_7_LFInst_0_n6,
         Red_PlaintextInst_LFInst_7_LFInst_0_n5,
         Red_PlaintextInst_LFInst_8_LFInst_0_n6,
         Red_PlaintextInst_LFInst_8_LFInst_0_n5,
         Red_PlaintextInst_LFInst_9_LFInst_0_n6,
         Red_PlaintextInst_LFInst_9_LFInst_0_n5,
         Red_PlaintextInst_LFInst_10_LFInst_0_n6,
         Red_PlaintextInst_LFInst_10_LFInst_0_n5,
         Red_PlaintextInst_LFInst_11_LFInst_0_n6,
         Red_PlaintextInst_LFInst_11_LFInst_0_n5,
         Red_PlaintextInst_LFInst_12_LFInst_0_n6,
         Red_PlaintextInst_LFInst_12_LFInst_0_n5,
         Red_PlaintextInst_LFInst_13_LFInst_0_n6,
         Red_PlaintextInst_LFInst_13_LFInst_0_n5,
         Red_PlaintextInst_LFInst_14_LFInst_0_n6,
         Red_PlaintextInst_LFInst_14_LFInst_0_n5,
         Red_PlaintextInst_LFInst_15_LFInst_0_n6,
         Red_PlaintextInst_LFInst_15_LFInst_0_n5,
         Red_SubCellInst_LFInst_0_LFInst_0_n9,
         Red_SubCellInst_LFInst_0_LFInst_0_n8,
         Red_SubCellInst_LFInst_0_LFInst_0_n7,
         Red_SubCellInst_LFInst_1_LFInst_0_n9,
         Red_SubCellInst_LFInst_1_LFInst_0_n8,
         Red_SubCellInst_LFInst_1_LFInst_0_n7,
         Red_SubCellInst_LFInst_2_LFInst_0_n9,
         Red_SubCellInst_LFInst_2_LFInst_0_n8,
         Red_SubCellInst_LFInst_2_LFInst_0_n7,
         Red_SubCellInst_LFInst_3_LFInst_0_n9,
         Red_SubCellInst_LFInst_3_LFInst_0_n8,
         Red_SubCellInst_LFInst_3_LFInst_0_n7,
         Red_SubCellInst_LFInst_4_LFInst_0_n9,
         Red_SubCellInst_LFInst_4_LFInst_0_n8,
         Red_SubCellInst_LFInst_4_LFInst_0_n7,
         Red_SubCellInst_LFInst_5_LFInst_0_n9,
         Red_SubCellInst_LFInst_5_LFInst_0_n8,
         Red_SubCellInst_LFInst_5_LFInst_0_n7,
         Red_SubCellInst_LFInst_6_LFInst_0_n9,
         Red_SubCellInst_LFInst_6_LFInst_0_n8,
         Red_SubCellInst_LFInst_6_LFInst_0_n7,
         Red_SubCellInst_LFInst_7_LFInst_0_n9,
         Red_SubCellInst_LFInst_7_LFInst_0_n8,
         Red_SubCellInst_LFInst_7_LFInst_0_n7,
         Red_SubCellInst_LFInst_8_LFInst_0_n9,
         Red_SubCellInst_LFInst_8_LFInst_0_n8,
         Red_SubCellInst_LFInst_8_LFInst_0_n7,
         Red_SubCellInst_LFInst_9_LFInst_0_n9,
         Red_SubCellInst_LFInst_9_LFInst_0_n8,
         Red_SubCellInst_LFInst_9_LFInst_0_n7,
         Red_SubCellInst_LFInst_10_LFInst_0_n9,
         Red_SubCellInst_LFInst_10_LFInst_0_n8,
         Red_SubCellInst_LFInst_10_LFInst_0_n7,
         Red_SubCellInst_LFInst_11_LFInst_0_n9,
         Red_SubCellInst_LFInst_11_LFInst_0_n8,
         Red_SubCellInst_LFInst_11_LFInst_0_n7,
         Red_SubCellInst_LFInst_12_LFInst_0_n9,
         Red_SubCellInst_LFInst_12_LFInst_0_n8,
         Red_SubCellInst_LFInst_12_LFInst_0_n7,
         Red_SubCellInst_LFInst_13_LFInst_0_n9,
         Red_SubCellInst_LFInst_13_LFInst_0_n8,
         Red_SubCellInst_LFInst_13_LFInst_0_n7,
         Red_SubCellInst_LFInst_14_LFInst_0_n9,
         Red_SubCellInst_LFInst_14_LFInst_0_n8,
         Red_SubCellInst_LFInst_14_LFInst_0_n7,
         Red_SubCellInst_LFInst_15_LFInst_0_n9,
         Red_SubCellInst_LFInst_15_LFInst_0_n8,
         Red_SubCellInst_LFInst_15_LFInst_0_n7, Red_MCInst_MC0_v3_3_0_,
         Red_MCInst_MC0_v3_2_0_, Red_MCInst_MC0_v3_1_0_,
         Red_MCInst_MC0_v3_0_0_, Red_MCInst_MC0_v2_3_0_,
         Red_MCInst_MC0_v2_2_0_, Red_MCInst_MC0_v2_1_0_,
         Red_MCInst_MC0_v2_0_0_, Red_MCInst_MC0_v1_3_0_,
         Red_MCInst_MC0_v1_2_0_, Red_MCInst_MC0_v1_1_0_,
         Red_MCInst_MC0_v1_0_0_, Red_MCInst_MC0_v0_3_0_,
         Red_MCInst_MC0_v0_2_0_, Red_MCInst_MC0_v0_1_0_,
         Red_MCInst_MC0_v0_0_0_, Red_MCInst_MC0_v0_3Inst_0_n3,
         Red_MCInst_MC0_v1_0Inst_0_n6, Red_MCInst_MC0_v1_0Inst_0_n5,
         Red_MCInst_MC0_v1_3Inst_0_n3, Red_MCInst_MC0_v2_0Inst_0_n3,
         Red_MCInst_MC0_v3_0Inst_0_n3, Red_MCInst_MC0_v3_2Inst_0_n3,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n7, Red_MCInst_MC1_v3_3_0_,
         Red_MCInst_MC1_v3_2_0_, Red_MCInst_MC1_v3_1_0_,
         Red_MCInst_MC1_v3_0_0_, Red_MCInst_MC1_v2_3_0_,
         Red_MCInst_MC1_v2_2_0_, Red_MCInst_MC1_v2_1_0_,
         Red_MCInst_MC1_v2_0_0_, Red_MCInst_MC1_v1_3_0_,
         Red_MCInst_MC1_v1_2_0_, Red_MCInst_MC1_v1_1_0_,
         Red_MCInst_MC1_v1_0_0_, Red_MCInst_MC1_v0_3_0_,
         Red_MCInst_MC1_v0_2_0_, Red_MCInst_MC1_v0_1_0_,
         Red_MCInst_MC1_v0_0_0_, Red_MCInst_MC1_v0_3Inst_0_n3,
         Red_MCInst_MC1_v1_0Inst_0_n6, Red_MCInst_MC1_v1_0Inst_0_n5,
         Red_MCInst_MC1_v1_3Inst_0_n3, Red_MCInst_MC1_v2_0Inst_0_n3,
         Red_MCInst_MC1_v3_0Inst_0_n3, Red_MCInst_MC1_v3_2Inst_0_n3,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n7, Red_MCInst_MC2_v3_3_0_,
         Red_MCInst_MC2_v3_2_0_, Red_MCInst_MC2_v3_1_0_,
         Red_MCInst_MC2_v3_0_0_, Red_MCInst_MC2_v2_3_0_,
         Red_MCInst_MC2_v2_2_0_, Red_MCInst_MC2_v2_1_0_,
         Red_MCInst_MC2_v2_0_0_, Red_MCInst_MC2_v1_3_0_,
         Red_MCInst_MC2_v1_2_0_, Red_MCInst_MC2_v1_1_0_,
         Red_MCInst_MC2_v1_0_0_, Red_MCInst_MC2_v0_3_0_,
         Red_MCInst_MC2_v0_2_0_, Red_MCInst_MC2_v0_1_0_,
         Red_MCInst_MC2_v0_0_0_, Red_MCInst_MC2_v0_3Inst_0_n3,
         Red_MCInst_MC2_v1_0Inst_0_n6, Red_MCInst_MC2_v1_0Inst_0_n5,
         Red_MCInst_MC2_v1_3Inst_0_n3, Red_MCInst_MC2_v2_0Inst_0_n3,
         Red_MCInst_MC2_v3_0Inst_0_n3, Red_MCInst_MC2_v3_2Inst_0_n3,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n7, Red_MCInst_MC3_v3_3_0_,
         Red_MCInst_MC3_v3_2_0_, Red_MCInst_MC3_v3_1_0_,
         Red_MCInst_MC3_v3_0_0_, Red_MCInst_MC3_v2_3_0_,
         Red_MCInst_MC3_v2_2_0_, Red_MCInst_MC3_v2_1_0_,
         Red_MCInst_MC3_v2_0_0_, Red_MCInst_MC3_v1_3_0_,
         Red_MCInst_MC3_v1_2_0_, Red_MCInst_MC3_v1_1_0_,
         Red_MCInst_MC3_v1_0_0_, Red_MCInst_MC3_v0_3_0_,
         Red_MCInst_MC3_v0_2_0_, Red_MCInst_MC3_v0_1_0_,
         Red_MCInst_MC3_v0_0_0_, Red_MCInst_MC3_v0_3Inst_0_n3,
         Red_MCInst_MC3_v1_0Inst_0_n6, Red_MCInst_MC3_v1_0Inst_0_n5,
         Red_MCInst_MC3_v1_3Inst_0_n3, Red_MCInst_MC3_v2_0Inst_0_n3,
         Red_MCInst_MC3_v3_0Inst_0_n3, Red_MCInst_MC3_v3_2Inst_0_n3,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n7,
         Red_SubCellInst2_LFInst_0_LFInst_0_n9,
         Red_SubCellInst2_LFInst_0_LFInst_0_n8,
         Red_SubCellInst2_LFInst_0_LFInst_0_n7,
         Red_SubCellInst2_LFInst_1_LFInst_0_n9,
         Red_SubCellInst2_LFInst_1_LFInst_0_n8,
         Red_SubCellInst2_LFInst_1_LFInst_0_n7,
         Red_SubCellInst2_LFInst_2_LFInst_0_n9,
         Red_SubCellInst2_LFInst_2_LFInst_0_n8,
         Red_SubCellInst2_LFInst_2_LFInst_0_n7,
         Red_SubCellInst2_LFInst_3_LFInst_0_n9,
         Red_SubCellInst2_LFInst_3_LFInst_0_n8,
         Red_SubCellInst2_LFInst_3_LFInst_0_n7,
         Red_SubCellInst2_LFInst_4_LFInst_0_n9,
         Red_SubCellInst2_LFInst_4_LFInst_0_n8,
         Red_SubCellInst2_LFInst_4_LFInst_0_n7,
         Red_SubCellInst2_LFInst_5_LFInst_0_n9,
         Red_SubCellInst2_LFInst_5_LFInst_0_n8,
         Red_SubCellInst2_LFInst_5_LFInst_0_n7,
         Red_SubCellInst2_LFInst_6_LFInst_0_n9,
         Red_SubCellInst2_LFInst_6_LFInst_0_n8,
         Red_SubCellInst2_LFInst_6_LFInst_0_n7,
         Red_SubCellInst2_LFInst_7_LFInst_0_n9,
         Red_SubCellInst2_LFInst_7_LFInst_0_n8,
         Red_SubCellInst2_LFInst_7_LFInst_0_n7,
         Red_SubCellInst2_LFInst_8_LFInst_0_n9,
         Red_SubCellInst2_LFInst_8_LFInst_0_n8,
         Red_SubCellInst2_LFInst_8_LFInst_0_n7,
         Red_SubCellInst2_LFInst_9_LFInst_0_n9,
         Red_SubCellInst2_LFInst_9_LFInst_0_n8,
         Red_SubCellInst2_LFInst_9_LFInst_0_n7,
         Red_SubCellInst2_LFInst_10_LFInst_0_n9,
         Red_SubCellInst2_LFInst_10_LFInst_0_n8,
         Red_SubCellInst2_LFInst_10_LFInst_0_n7,
         Red_SubCellInst2_LFInst_11_LFInst_0_n9,
         Red_SubCellInst2_LFInst_11_LFInst_0_n8,
         Red_SubCellInst2_LFInst_11_LFInst_0_n7,
         Red_SubCellInst2_LFInst_12_LFInst_0_n9,
         Red_SubCellInst2_LFInst_12_LFInst_0_n8,
         Red_SubCellInst2_LFInst_12_LFInst_0_n7,
         Red_SubCellInst2_LFInst_13_LFInst_0_n9,
         Red_SubCellInst2_LFInst_13_LFInst_0_n8,
         Red_SubCellInst2_LFInst_13_LFInst_0_n7,
         Red_SubCellInst2_LFInst_14_LFInst_0_n9,
         Red_SubCellInst2_LFInst_14_LFInst_0_n8,
         Red_SubCellInst2_LFInst_14_LFInst_0_n7,
         Red_SubCellInst2_LFInst_15_LFInst_0_n9,
         Red_SubCellInst2_LFInst_15_LFInst_0_n8,
         Red_SubCellInst2_LFInst_15_LFInst_0_n7, Red_MCInst2_MC0_v3_3_0_,
         Red_MCInst2_MC0_v3_2_0_, Red_MCInst2_MC0_v3_1_0_,
         Red_MCInst2_MC0_v3_0_0_, Red_MCInst2_MC0_v2_3_0_,
         Red_MCInst2_MC0_v2_2_0_, Red_MCInst2_MC0_v2_1_0_,
         Red_MCInst2_MC0_v2_0_0_, Red_MCInst2_MC0_v1_3_0_,
         Red_MCInst2_MC0_v1_2_0_, Red_MCInst2_MC0_v1_1_0_,
         Red_MCInst2_MC0_v1_0_0_, Red_MCInst2_MC0_v0_3_0_,
         Red_MCInst2_MC0_v0_2_0_, Red_MCInst2_MC0_v0_1_0_,
         Red_MCInst2_MC0_v0_0_0_, Red_MCInst2_MC0_v0_3Inst_0_n3,
         Red_MCInst2_MC0_v1_0Inst_0_n6, Red_MCInst2_MC0_v1_0Inst_0_n5,
         Red_MCInst2_MC0_v1_3Inst_0_n3, Red_MCInst2_MC0_v2_0Inst_0_n3,
         Red_MCInst2_MC0_v3_0Inst_0_n3, Red_MCInst2_MC0_v3_2Inst_0_n3,
         Red_MCInst2_MC0_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r3Inst_XORInst_0_0_n7, Red_MCInst2_MC1_v3_3_0_,
         Red_MCInst2_MC1_v3_2_0_, Red_MCInst2_MC1_v3_1_0_,
         Red_MCInst2_MC1_v3_0_0_, Red_MCInst2_MC1_v2_3_0_,
         Red_MCInst2_MC1_v2_2_0_, Red_MCInst2_MC1_v2_1_0_,
         Red_MCInst2_MC1_v2_0_0_, Red_MCInst2_MC1_v1_3_0_,
         Red_MCInst2_MC1_v1_2_0_, Red_MCInst2_MC1_v1_1_0_,
         Red_MCInst2_MC1_v1_0_0_, Red_MCInst2_MC1_v0_3_0_,
         Red_MCInst2_MC1_v0_2_0_, Red_MCInst2_MC1_v0_1_0_,
         Red_MCInst2_MC1_v0_0_0_, Red_MCInst2_MC1_v0_3Inst_0_n3,
         Red_MCInst2_MC1_v1_0Inst_0_n6, Red_MCInst2_MC1_v1_0Inst_0_n5,
         Red_MCInst2_MC1_v1_3Inst_0_n3, Red_MCInst2_MC1_v2_0Inst_0_n3,
         Red_MCInst2_MC1_v3_0Inst_0_n3, Red_MCInst2_MC1_v3_2Inst_0_n3,
         Red_MCInst2_MC1_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r3Inst_XORInst_0_0_n7, Red_MCInst2_MC2_v3_3_0_,
         Red_MCInst2_MC2_v3_2_0_, Red_MCInst2_MC2_v3_1_0_,
         Red_MCInst2_MC2_v3_0_0_, Red_MCInst2_MC2_v2_3_0_,
         Red_MCInst2_MC2_v2_2_0_, Red_MCInst2_MC2_v2_1_0_,
         Red_MCInst2_MC2_v2_0_0_, Red_MCInst2_MC2_v1_3_0_,
         Red_MCInst2_MC2_v1_2_0_, Red_MCInst2_MC2_v1_1_0_,
         Red_MCInst2_MC2_v1_0_0_, Red_MCInst2_MC2_v0_3_0_,
         Red_MCInst2_MC2_v0_2_0_, Red_MCInst2_MC2_v0_1_0_,
         Red_MCInst2_MC2_v0_0_0_, Red_MCInst2_MC2_v0_3Inst_0_n3,
         Red_MCInst2_MC2_v1_0Inst_0_n6, Red_MCInst2_MC2_v1_0Inst_0_n5,
         Red_MCInst2_MC2_v1_3Inst_0_n3, Red_MCInst2_MC2_v2_0Inst_0_n3,
         Red_MCInst2_MC2_v3_0Inst_0_n3, Red_MCInst2_MC2_v3_2Inst_0_n3,
         Red_MCInst2_MC2_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r3Inst_XORInst_0_0_n7, Red_MCInst2_MC3_v3_3_0_,
         Red_MCInst2_MC3_v3_2_0_, Red_MCInst2_MC3_v3_1_0_,
         Red_MCInst2_MC3_v3_0_0_, Red_MCInst2_MC3_v2_3_0_,
         Red_MCInst2_MC3_v2_2_0_, Red_MCInst2_MC3_v2_1_0_,
         Red_MCInst2_MC3_v2_0_0_, Red_MCInst2_MC3_v1_3_0_,
         Red_MCInst2_MC3_v1_2_0_, Red_MCInst2_MC3_v1_1_0_,
         Red_MCInst2_MC3_v1_0_0_, Red_MCInst2_MC3_v0_3_0_,
         Red_MCInst2_MC3_v0_2_0_, Red_MCInst2_MC3_v0_1_0_,
         Red_MCInst2_MC3_v0_0_0_, Red_MCInst2_MC3_v0_3Inst_0_n3,
         Red_MCInst2_MC3_v1_0Inst_0_n6, Red_MCInst2_MC3_v1_0Inst_0_n5,
         Red_MCInst2_MC3_v1_3Inst_0_n3, Red_MCInst2_MC3_v2_0Inst_0_n3,
         Red_MCInst2_MC3_v3_0Inst_0_n3, Red_MCInst2_MC3_v3_2Inst_0_n3,
         Red_MCInst2_MC3_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r3Inst_XORInst_0_0_n7,
         Red_KeyInst_LFInst_0_LFInst_0_n6, Red_KeyInst_LFInst_0_LFInst_0_n5,
         Red_KeyInst_LFInst_1_LFInst_0_n6, Red_KeyInst_LFInst_1_LFInst_0_n5,
         Red_KeyInst_LFInst_2_LFInst_0_n6, Red_KeyInst_LFInst_2_LFInst_0_n5,
         Red_KeyInst_LFInst_3_LFInst_0_n6, Red_KeyInst_LFInst_3_LFInst_0_n5,
         Red_KeyInst_LFInst_4_LFInst_0_n6, Red_KeyInst_LFInst_4_LFInst_0_n5,
         Red_KeyInst_LFInst_5_LFInst_0_n6, Red_KeyInst_LFInst_5_LFInst_0_n5,
         Red_KeyInst_LFInst_6_LFInst_0_n6, Red_KeyInst_LFInst_6_LFInst_0_n5,
         Red_KeyInst_LFInst_7_LFInst_0_n6, Red_KeyInst_LFInst_7_LFInst_0_n5,
         Red_KeyInst_LFInst_8_LFInst_0_n6, Red_KeyInst_LFInst_8_LFInst_0_n5,
         Red_KeyInst_LFInst_9_LFInst_0_n6, Red_KeyInst_LFInst_9_LFInst_0_n5,
         Red_KeyInst_LFInst_10_LFInst_0_n6, Red_KeyInst_LFInst_10_LFInst_0_n5,
         Red_KeyInst_LFInst_11_LFInst_0_n6, Red_KeyInst_LFInst_11_LFInst_0_n5,
         Red_KeyInst_LFInst_12_LFInst_0_n6, Red_KeyInst_LFInst_12_LFInst_0_n5,
         Red_KeyInst_LFInst_13_LFInst_0_n6, Red_KeyInst_LFInst_13_LFInst_0_n5,
         Red_KeyInst_LFInst_14_LFInst_0_n6, Red_KeyInst_LFInst_14_LFInst_0_n5,
         Red_KeyInst_LFInst_15_LFInst_0_n6, Red_KeyInst_LFInst_15_LFInst_0_n5,
         Red_ToCheckInst_LFInst_0_LFInst_0_n6,
         Red_ToCheckInst_LFInst_0_LFInst_0_n5,
         Red_ToCheckInst_LFInst_1_LFInst_0_n6,
         Red_ToCheckInst_LFInst_1_LFInst_0_n5,
         Red_ToCheckInst_LFInst_2_LFInst_0_n6,
         Red_ToCheckInst_LFInst_2_LFInst_0_n5,
         Red_ToCheckInst_LFInst_3_LFInst_0_n6,
         Red_ToCheckInst_LFInst_3_LFInst_0_n5,
         Red_ToCheckInst_LFInst_4_LFInst_0_n6,
         Red_ToCheckInst_LFInst_4_LFInst_0_n5,
         Red_ToCheckInst_LFInst_5_LFInst_0_n6,
         Red_ToCheckInst_LFInst_5_LFInst_0_n5,
         Red_ToCheckInst_LFInst_6_LFInst_0_n6,
         Red_ToCheckInst_LFInst_6_LFInst_0_n5,
         Red_ToCheckInst_LFInst_7_LFInst_0_n6,
         Red_ToCheckInst_LFInst_7_LFInst_0_n5,
         Red_ToCheckInst_LFInst_8_LFInst_0_n6,
         Red_ToCheckInst_LFInst_8_LFInst_0_n5,
         Red_ToCheckInst_LFInst_9_LFInst_0_n6,
         Red_ToCheckInst_LFInst_9_LFInst_0_n5,
         Red_ToCheckInst_LFInst_10_LFInst_0_n6,
         Red_ToCheckInst_LFInst_10_LFInst_0_n5,
         Red_ToCheckInst_LFInst_11_LFInst_0_n6,
         Red_ToCheckInst_LFInst_11_LFInst_0_n5,
         Red_ToCheckInst_LFInst_12_LFInst_0_n6,
         Red_ToCheckInst_LFInst_12_LFInst_0_n5,
         Red_ToCheckInst_LFInst_13_LFInst_0_n6,
         Red_ToCheckInst_LFInst_13_LFInst_0_n5,
         Red_ToCheckInst_LFInst_14_LFInst_0_n6,
         Red_ToCheckInst_LFInst_14_LFInst_0_n5,
         Red_ToCheckInst_LFInst_15_LFInst_0_n6,
         Red_ToCheckInst_LFInst_15_LFInst_0_n5,
         Red_ToCheckInst_LFInst_16_LFInst_0_n6,
         Red_ToCheckInst_LFInst_16_LFInst_0_n5,
         Red_ToCheckInst_LFInst_17_LFInst_0_n6,
         Red_ToCheckInst_LFInst_17_LFInst_0_n5,
         Red_ToCheckInst_LFInst_18_LFInst_0_n6,
         Red_ToCheckInst_LFInst_18_LFInst_0_n5,
         Red_ToCheckInst_LFInst_19_LFInst_0_n6,
         Red_ToCheckInst_LFInst_19_LFInst_0_n5,
         Red_ToCheckInst_LFInst_20_LFInst_0_n6,
         Red_ToCheckInst_LFInst_20_LFInst_0_n5,
         Red_ToCheckInst_LFInst_21_LFInst_0_n6,
         Red_ToCheckInst_LFInst_21_LFInst_0_n5,
         Red_ToCheckInst_LFInst_22_LFInst_0_n6,
         Red_ToCheckInst_LFInst_22_LFInst_0_n5,
         Red_ToCheckInst_LFInst_23_LFInst_0_n6,
         Red_ToCheckInst_LFInst_23_LFInst_0_n5,
         Red_ToCheckInst_LFInst_24_LFInst_0_n6,
         Red_ToCheckInst_LFInst_24_LFInst_0_n5,
         Red_ToCheckInst_LFInst_25_LFInst_0_n6,
         Red_ToCheckInst_LFInst_25_LFInst_0_n5,
         Red_ToCheckInst_LFInst_26_LFInst_0_n6,
         Red_ToCheckInst_LFInst_26_LFInst_0_n5,
         Red_ToCheckInst_LFInst_27_LFInst_0_n6,
         Red_ToCheckInst_LFInst_27_LFInst_0_n5,
         Red_ToCheckInst_LFInst_28_LFInst_0_n6,
         Red_ToCheckInst_LFInst_28_LFInst_0_n5,
         Red_ToCheckInst_LFInst_29_LFInst_0_n6,
         Red_ToCheckInst_LFInst_29_LFInst_0_n5,
         Red_ToCheckInst_LFInst_30_LFInst_0_n6,
         Red_ToCheckInst_LFInst_30_LFInst_0_n5,
         Red_ToCheckInst_LFInst_31_LFInst_0_n6,
         Red_ToCheckInst_LFInst_31_LFInst_0_n5,
         Red_ToCheckInst_LFInst_32_LFInst_0_n6,
         Red_ToCheckInst_LFInst_32_LFInst_0_n5,
         Red_ToCheckInst_LFInst_33_LFInst_0_n6,
         Red_ToCheckInst_LFInst_33_LFInst_0_n5,
         Red_ToCheckInst_LFInst_34_LFInst_0_n6,
         Red_ToCheckInst_LFInst_34_LFInst_0_n5,
         Red_ToCheckInst_LFInst_35_LFInst_0_n6,
         Red_ToCheckInst_LFInst_35_LFInst_0_n5,
         Red_ToCheckInst_LFInst_36_LFInst_0_n6,
         Red_ToCheckInst_LFInst_36_LFInst_0_n5,
         Red_ToCheckInst_LFInst_37_LFInst_0_n6,
         Red_ToCheckInst_LFInst_37_LFInst_0_n5,
         Red_ToCheckInst_LFInst_38_LFInst_0_n6,
         Red_ToCheckInst_LFInst_38_LFInst_0_n5,
         Red_ToCheckInst_LFInst_39_LFInst_0_n6,
         Red_ToCheckInst_LFInst_39_LFInst_0_n5,
         Red_ToCheckInst_LFInst_40_LFInst_0_n6,
         Red_ToCheckInst_LFInst_40_LFInst_0_n5,
         Red_ToCheckInst_LFInst_41_LFInst_0_n6,
         Red_ToCheckInst_LFInst_41_LFInst_0_n5,
         Red_ToCheckInst_LFInst_42_LFInst_0_n6,
         Red_ToCheckInst_LFInst_42_LFInst_0_n5,
         Red_ToCheckInst_LFInst_43_LFInst_0_n6,
         Red_ToCheckInst_LFInst_43_LFInst_0_n5,
         Red_ToCheckInst_LFInst_44_LFInst_0_n6,
         Red_ToCheckInst_LFInst_44_LFInst_0_n5,
         Red_ToCheckInst_LFInst_45_LFInst_0_n6,
         Red_ToCheckInst_LFInst_45_LFInst_0_n5,
         Red_ToCheckInst_LFInst_46_LFInst_0_n6,
         Red_ToCheckInst_LFInst_46_LFInst_0_n5,
         Red_ToCheckInst_LFInst_47_LFInst_0_n6,
         Red_ToCheckInst_LFInst_47_LFInst_0_n5,
         Red_ToCheckInst_LFInst_48_LFInst_0_n6,
         Red_ToCheckInst_LFInst_48_LFInst_0_n5,
         Red_ToCheckInst_LFInst_49_LFInst_0_n6,
         Red_ToCheckInst_LFInst_49_LFInst_0_n5,
         Red_ToCheckInst_LFInst_50_LFInst_0_n6,
         Red_ToCheckInst_LFInst_50_LFInst_0_n5,
         Red_ToCheckInst_LFInst_51_LFInst_0_n6,
         Red_ToCheckInst_LFInst_51_LFInst_0_n5,
         Red_ToCheckInst_LFInst_52_LFInst_0_n6,
         Red_ToCheckInst_LFInst_52_LFInst_0_n5,
         Red_ToCheckInst_LFInst_53_LFInst_0_n6,
         Red_ToCheckInst_LFInst_53_LFInst_0_n5,
         Red_ToCheckInst_LFInst_54_LFInst_0_n6,
         Red_ToCheckInst_LFInst_54_LFInst_0_n5,
         Red_ToCheckInst_LFInst_55_LFInst_0_n6,
         Red_ToCheckInst_LFInst_55_LFInst_0_n5,
         Red_ToCheckInst_LFInst_56_LFInst_0_n6,
         Red_ToCheckInst_LFInst_56_LFInst_0_n5,
         Red_ToCheckInst_LFInst_57_LFInst_0_n6,
         Red_ToCheckInst_LFInst_57_LFInst_0_n5,
         Red_ToCheckInst_LFInst_58_LFInst_0_n6,
         Red_ToCheckInst_LFInst_58_LFInst_0_n5,
         Red_ToCheckInst_LFInst_59_LFInst_0_n6,
         Red_ToCheckInst_LFInst_59_LFInst_0_n5,
         Red_ToCheckInst_LFInst_60_LFInst_0_n6,
         Red_ToCheckInst_LFInst_60_LFInst_0_n5,
         Red_ToCheckInst_LFInst_61_LFInst_0_n6,
         Red_ToCheckInst_LFInst_61_LFInst_0_n5,
         Red_ToCheckInst_LFInst_62_LFInst_0_n6,
         Red_ToCheckInst_LFInst_62_LFInst_0_n5,
         Red_ToCheckInst_LFInst_63_LFInst_0_n6,
         Red_ToCheckInst_LFInst_63_LFInst_0_n5,
         Red_ToCheckInst_LFInst_64_LFInst_0_n6,
         Red_ToCheckInst_LFInst_64_LFInst_0_n5,
         Red_ToCheckInst_LFInst_65_LFInst_0_n6,
         Red_ToCheckInst_LFInst_65_LFInst_0_n5,
         Red_ToCheckInst_LFInst_66_LFInst_0_n6,
         Red_ToCheckInst_LFInst_66_LFInst_0_n5,
         Red_ToCheckInst_LFInst_67_LFInst_0_n6,
         Red_ToCheckInst_LFInst_67_LFInst_0_n5,
         Red_ToCheckInst_LFInst_68_LFInst_0_n6,
         Red_ToCheckInst_LFInst_68_LFInst_0_n5,
         Red_ToCheckInst_LFInst_69_LFInst_0_n6,
         Red_ToCheckInst_LFInst_69_LFInst_0_n5,
         Red_ToCheckInst_LFInst_70_LFInst_0_n6,
         Red_ToCheckInst_LFInst_70_LFInst_0_n5,
         Red_ToCheckInst_LFInst_71_LFInst_0_n6,
         Red_ToCheckInst_LFInst_71_LFInst_0_n5,
         Red_ToCheckInst_LFInst_72_LFInst_0_n6,
         Red_ToCheckInst_LFInst_72_LFInst_0_n5,
         Red_ToCheckInst_LFInst_73_LFInst_0_n6,
         Red_ToCheckInst_LFInst_73_LFInst_0_n5,
         Red_ToCheckInst_LFInst_74_LFInst_0_n6,
         Red_ToCheckInst_LFInst_74_LFInst_0_n5,
         Red_ToCheckInst_LFInst_75_LFInst_0_n6,
         Red_ToCheckInst_LFInst_75_LFInst_0_n5,
         Red_ToCheckInst_LFInst_76_LFInst_0_n6,
         Red_ToCheckInst_LFInst_76_LFInst_0_n5,
         Red_ToCheckInst_LFInst_77_LFInst_0_n6,
         Red_ToCheckInst_LFInst_77_LFInst_0_n5,
         Red_ToCheckInst_LFInst_78_LFInst_0_n6,
         Red_ToCheckInst_LFInst_78_LFInst_0_n5,
         Red_ToCheckInst_LFInst_79_LFInst_0_n6,
         Red_ToCheckInst_LFInst_79_LFInst_0_n5,
         Red_ToCheckInst_LFInst_80_LFInst_0_n6,
         Red_ToCheckInst_LFInst_80_LFInst_0_n5,
         Red_ToCheckInst_LFInst_81_LFInst_0_n6,
         Red_ToCheckInst_LFInst_81_LFInst_0_n5,
         Red_ToCheckInst_LFInst_82_LFInst_0_n6,
         Red_ToCheckInst_LFInst_82_LFInst_0_n5,
         Red_ToCheckInst_LFInst_83_LFInst_0_n6,
         Red_ToCheckInst_LFInst_83_LFInst_0_n5,
         Red_ToCheckInst_LFInst_84_LFInst_0_n6,
         Red_ToCheckInst_LFInst_84_LFInst_0_n5,
         Red_ToCheckInst_LFInst_85_LFInst_0_n6,
         Red_ToCheckInst_LFInst_85_LFInst_0_n5,
         Red_ToCheckInst_LFInst_86_LFInst_0_n6,
         Red_ToCheckInst_LFInst_86_LFInst_0_n5,
         Red_ToCheckInst_LFInst_87_LFInst_0_n6,
         Red_ToCheckInst_LFInst_87_LFInst_0_n5,
         Red_ToCheckInst_LFInst_88_LFInst_0_n6,
         Red_ToCheckInst_LFInst_88_LFInst_0_n5,
         Red_ToCheckInst_LFInst_89_LFInst_0_n6,
         Red_ToCheckInst_LFInst_89_LFInst_0_n5,
         Red_ToCheckInst_LFInst_90_LFInst_0_n6,
         Red_ToCheckInst_LFInst_90_LFInst_0_n5,
         Red_ToCheckInst_LFInst_91_LFInst_0_n6,
         Red_ToCheckInst_LFInst_91_LFInst_0_n5,
         Red_ToCheckInst_LFInst_92_LFInst_0_n6,
         Red_ToCheckInst_LFInst_92_LFInst_0_n5,
         Red_ToCheckInst_LFInst_93_LFInst_0_n6,
         Red_ToCheckInst_LFInst_93_LFInst_0_n5,
         Red_ToCheckInst_LFInst_94_LFInst_0_n6,
         Red_ToCheckInst_LFInst_94_LFInst_0_n5,
         Red_ToCheckInst_LFInst_95_LFInst_0_n6,
         Red_ToCheckInst_LFInst_95_LFInst_0_n5, Check1_CheckInst_0_n190,
         Check1_CheckInst_0_n189, Check1_CheckInst_0_n188,
         Check1_CheckInst_0_n187, Check1_CheckInst_0_n186,
         Check1_CheckInst_0_n185, Check1_CheckInst_0_n184,
         Check1_CheckInst_0_n183, Check1_CheckInst_0_n182,
         Check1_CheckInst_0_n181, Check1_CheckInst_0_n180,
         Check1_CheckInst_0_n179, Check1_CheckInst_0_n178,
         Check1_CheckInst_0_n177, Check1_CheckInst_0_n176,
         Check1_CheckInst_0_n175, Check1_CheckInst_0_n174,
         Check1_CheckInst_0_n173, Check1_CheckInst_0_n172,
         Check1_CheckInst_0_n171, Check1_CheckInst_0_n170,
         Check1_CheckInst_0_n169, Check1_CheckInst_0_n168,
         Check1_CheckInst_0_n167, Check1_CheckInst_0_n166,
         Check1_CheckInst_0_n165, Check1_CheckInst_0_n164,
         Check1_CheckInst_0_n163, Check1_CheckInst_0_n162,
         Check1_CheckInst_0_n161, Check1_CheckInst_0_n160,
         Check1_CheckInst_0_n159, Check1_CheckInst_0_n158,
         Check1_CheckInst_0_n157, Check1_CheckInst_0_n156,
         Check1_CheckInst_0_n155, Check1_CheckInst_0_n154,
         Check1_CheckInst_0_n153, Check1_CheckInst_0_n152,
         Check1_CheckInst_0_n151, Check1_CheckInst_0_n150,
         Check1_CheckInst_0_n149, Check1_CheckInst_0_n148,
         Check1_CheckInst_0_n147, Check1_CheckInst_0_n146,
         Check1_CheckInst_0_n145, Check1_CheckInst_0_n144,
         Check1_CheckInst_0_n143, Check1_CheckInst_0_n142,
         Check1_CheckInst_0_n141, Check1_CheckInst_0_n140,
         Check1_CheckInst_0_n139, Check1_CheckInst_0_n138,
         Check1_CheckInst_0_n137, Check1_CheckInst_0_n136,
         Check1_CheckInst_0_n135, Check1_CheckInst_0_n134,
         Check1_CheckInst_0_n133, Check1_CheckInst_0_n132,
         Check1_CheckInst_0_n131, Check1_CheckInst_0_n130,
         Check1_CheckInst_0_n129, Check1_CheckInst_0_n128,
         Check1_CheckInst_0_n127, Check1_CheckInst_0_n126,
         Check1_CheckInst_0_n125, Check1_CheckInst_0_n124,
         Check1_CheckInst_0_n123, Check1_CheckInst_0_n122,
         Check1_CheckInst_0_n121, Check1_CheckInst_0_n120,
         Check1_CheckInst_0_n119, Check1_CheckInst_0_n118,
         Check1_CheckInst_0_n117, Check1_CheckInst_0_n116,
         Check1_CheckInst_0_n115, Check1_CheckInst_0_n114,
         Check1_CheckInst_0_n113, Check1_CheckInst_0_n112,
         Check1_CheckInst_0_n111, Check1_CheckInst_0_n110,
         Check1_CheckInst_0_n109, Check1_CheckInst_0_n108,
         Check1_CheckInst_0_n107, Check1_CheckInst_0_n106,
         Check1_CheckInst_0_n105, Check1_CheckInst_0_n104,
         Check1_CheckInst_0_n103, Check1_CheckInst_0_n102,
         Check1_CheckInst_0_n101, Check1_CheckInst_0_n100,
         Check1_CheckInst_0_n99, Check1_CheckInst_0_n98,
         Check1_CheckInst_0_n97, Check1_CheckInst_0_n96,
         Check1_CheckInst_0_n95, Check1_CheckInst_0_n94,
         Check1_CheckInst_0_n93, Check1_CheckInst_0_n92,
         Check1_CheckInst_0_n91, Check1_CheckInst_0_n90,
         Check1_CheckInst_0_n89, Check1_CheckInst_0_n88,
         Check1_CheckInst_0_n87, Check1_CheckInst_0_n86,
         Check1_CheckInst_0_n85, Check1_CheckInst_0_n84,
         Check1_CheckInst_0_n83, Check1_CheckInst_0_n82,
         Check1_CheckInst_0_n81, Check1_CheckInst_0_n80,
         Check1_CheckInst_0_n79, Check1_CheckInst_0_n78,
         Check1_CheckInst_0_n77, Check1_CheckInst_0_n76,
         Check1_CheckInst_0_n75, Check1_CheckInst_0_n74,
         Check1_CheckInst_0_n73, Check1_CheckInst_0_n72,
         Check1_CheckInst_0_n71, Check1_CheckInst_0_n70,
         Check1_CheckInst_0_n69, Check1_CheckInst_0_n68,
         Check1_CheckInst_0_n67, Check1_CheckInst_0_n66,
         Check1_CheckInst_0_n65, Check1_CheckInst_0_n64,
         Check1_CheckInst_0_n63, Check1_CheckInst_0_n62,
         Check1_CheckInst_0_n61, Check1_CheckInst_0_n60,
         Check1_CheckInst_0_n59, Check1_CheckInst_0_n58,
         Check1_CheckInst_0_n57, Check1_CheckInst_0_n56,
         Check1_CheckInst_0_n55, Check1_CheckInst_0_n54,
         Check1_CheckInst_0_n53, Check1_CheckInst_0_n52,
         Check1_CheckInst_0_n51, Check1_CheckInst_0_n50,
         Check1_CheckInst_0_n49, Check1_CheckInst_0_n48,
         Check1_CheckInst_0_n47, Check1_CheckInst_0_n46,
         Check1_CheckInst_0_n45, Check1_CheckInst_0_n44,
         Check1_CheckInst_0_n43, Check1_CheckInst_0_n42,
         Check1_CheckInst_0_n41, Check1_CheckInst_0_n40,
         Check1_CheckInst_0_n39, Check1_CheckInst_0_n38,
         Check1_CheckInst_0_n37, Check1_CheckInst_0_n36,
         Check1_CheckInst_0_n35, Check1_CheckInst_0_n34,
         Check1_CheckInst_0_n33, Check1_CheckInst_0_n32,
         Check1_CheckInst_0_n31, Check1_CheckInst_0_n30,
         Check1_CheckInst_0_n29, Check1_CheckInst_0_n28,
         Check1_CheckInst_0_n27, Check1_CheckInst_0_n26,
         Check1_CheckInst_0_n25, Check1_CheckInst_0_n24,
         Check1_CheckInst_0_n23, Check1_CheckInst_0_n22,
         Check1_CheckInst_0_n21, Check1_CheckInst_0_n20,
         Check1_CheckInst_0_n19, Check1_CheckInst_0_n18,
         Check1_CheckInst_0_n17, Check1_CheckInst_0_n16,
         Check1_CheckInst_0_n15, Check1_CheckInst_0_n14,
         Check1_CheckInst_0_n13, Check1_CheckInst_0_n12,
         Check1_CheckInst_0_n11, Check1_CheckInst_0_n10, Check1_CheckInst_0_n9,
         Check1_CheckInst_0_n8, Check1_CheckInst_0_n7, Check1_CheckInst_0_n6,
         Check1_CheckInst_0_n5, Check1_CheckInst_0_n4, Check1_CheckInst_0_n3,
         Check1_CheckInst_0_n2, Check1_CheckInst_0_n1;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] MC_output;
  wire   [63:0] SubCellInput2;
  wire   [15:0] Red_Plaintext;
  wire   [15:0] Red_RoundKey;
  wire   [15:0] Red_AddRoundKeyOutput;
  wire   [15:0] Red_ShiftRowsOutput;
  wire   [15:0] Red_MC_output;
  wire   [15:0] Red_SubCellInput2;
  wire   [15:0] Red_ShiftRowsOutput2;
  wire   [15:0] Red_MC_output2;
  wire   [95:0] Red_SignaltoCheck;
  wire   [3:0] MCInst_MC0_v3_3;
  wire   [3:0] MCInst_MC0_v3_2;
  wire   [3:0] MCInst_MC0_v3_1;
  wire   [2:1] MCInst_MC0_v3_0;
  wire   [3:0] MCInst_MC0_v2_3;
  wire   [3:0] MCInst_MC0_v2_2;
  wire   [3:0] MCInst_MC0_v2_1;
  wire   [3:0] MCInst_MC0_v2_0;
  wire   [2:1] MCInst_MC0_v1_3;
  wire   [3:0] MCInst_MC0_v1_2;
  wire   [3:0] MCInst_MC0_v1_1;
  wire   [3:0] MCInst_MC0_v1_0;
  wire   [3:0] MCInst_MC0_v0_3;
  wire   [3:0] MCInst_MC0_v0_2;
  wire   [3:1] MCInst_MC0_v0_1;
  wire   [3:1] MCInst_MC0_v0_0;
  wire   [3:0] MCInst_MC1_v3_3;
  wire   [3:0] MCInst_MC1_v3_2;
  wire   [3:0] MCInst_MC1_v3_1;
  wire   [2:1] MCInst_MC1_v3_0;
  wire   [3:0] MCInst_MC1_v2_3;
  wire   [3:0] MCInst_MC1_v2_2;
  wire   [3:0] MCInst_MC1_v2_1;
  wire   [3:0] MCInst_MC1_v2_0;
  wire   [2:1] MCInst_MC1_v1_3;
  wire   [3:0] MCInst_MC1_v1_2;
  wire   [3:0] MCInst_MC1_v1_1;
  wire   [3:0] MCInst_MC1_v1_0;
  wire   [3:0] MCInst_MC1_v0_3;
  wire   [3:0] MCInst_MC1_v0_2;
  wire   [3:1] MCInst_MC1_v0_1;
  wire   [3:1] MCInst_MC1_v0_0;
  wire   [3:0] MCInst_MC2_v3_3;
  wire   [3:0] MCInst_MC2_v3_2;
  wire   [3:0] MCInst_MC2_v3_1;
  wire   [2:1] MCInst_MC2_v3_0;
  wire   [3:0] MCInst_MC2_v2_3;
  wire   [3:0] MCInst_MC2_v2_2;
  wire   [3:0] MCInst_MC2_v2_1;
  wire   [3:0] MCInst_MC2_v2_0;
  wire   [2:1] MCInst_MC2_v1_3;
  wire   [3:0] MCInst_MC2_v1_2;
  wire   [3:0] MCInst_MC2_v1_1;
  wire   [3:0] MCInst_MC2_v1_0;
  wire   [3:0] MCInst_MC2_v0_3;
  wire   [3:0] MCInst_MC2_v0_2;
  wire   [3:1] MCInst_MC2_v0_1;
  wire   [3:1] MCInst_MC2_v0_0;
  wire   [3:0] MCInst_MC3_v3_3;
  wire   [3:0] MCInst_MC3_v3_2;
  wire   [3:0] MCInst_MC3_v3_1;
  wire   [2:1] MCInst_MC3_v3_0;
  wire   [3:0] MCInst_MC3_v2_3;
  wire   [3:0] MCInst_MC3_v2_2;
  wire   [3:0] MCInst_MC3_v2_1;
  wire   [3:0] MCInst_MC3_v2_0;
  wire   [2:1] MCInst_MC3_v1_3;
  wire   [3:0] MCInst_MC3_v1_2;
  wire   [3:0] MCInst_MC3_v1_1;
  wire   [3:0] MCInst_MC3_v1_0;
  wire   [3:0] MCInst_MC3_v0_3;
  wire   [3:0] MCInst_MC3_v0_2;
  wire   [3:1] MCInst_MC3_v0_1;
  wire   [3:1] MCInst_MC3_v0_0;
  wire   [3:0] MCInst2_MC0_v3_3;
  wire   [3:0] MCInst2_MC0_v3_2;
  wire   [3:0] MCInst2_MC0_v3_1;
  wire   [2:1] MCInst2_MC0_v3_0;
  wire   [3:0] MCInst2_MC0_v2_3;
  wire   [3:0] MCInst2_MC0_v2_2;
  wire   [3:0] MCInst2_MC0_v2_1;
  wire   [3:0] MCInst2_MC0_v2_0;
  wire   [2:1] MCInst2_MC0_v1_3;
  wire   [3:0] MCInst2_MC0_v1_2;
  wire   [3:0] MCInst2_MC0_v1_1;
  wire   [3:0] MCInst2_MC0_v1_0;
  wire   [3:0] MCInst2_MC0_v0_3;
  wire   [3:0] MCInst2_MC0_v0_2;
  wire   [3:1] MCInst2_MC0_v0_1;
  wire   [3:1] MCInst2_MC0_v0_0;
  wire   [3:0] MCInst2_MC1_v3_3;
  wire   [3:0] MCInst2_MC1_v3_2;
  wire   [3:0] MCInst2_MC1_v3_1;
  wire   [2:1] MCInst2_MC1_v3_0;
  wire   [3:0] MCInst2_MC1_v2_3;
  wire   [3:0] MCInst2_MC1_v2_2;
  wire   [3:0] MCInst2_MC1_v2_1;
  wire   [3:0] MCInst2_MC1_v2_0;
  wire   [2:1] MCInst2_MC1_v1_3;
  wire   [3:0] MCInst2_MC1_v1_2;
  wire   [3:0] MCInst2_MC1_v1_1;
  wire   [3:0] MCInst2_MC1_v1_0;
  wire   [3:0] MCInst2_MC1_v0_3;
  wire   [3:0] MCInst2_MC1_v0_2;
  wire   [3:1] MCInst2_MC1_v0_1;
  wire   [3:1] MCInst2_MC1_v0_0;
  wire   [3:0] MCInst2_MC2_v3_3;
  wire   [3:0] MCInst2_MC2_v3_2;
  wire   [3:0] MCInst2_MC2_v3_1;
  wire   [2:1] MCInst2_MC2_v3_0;
  wire   [3:0] MCInst2_MC2_v2_3;
  wire   [3:0] MCInst2_MC2_v2_2;
  wire   [3:0] MCInst2_MC2_v2_1;
  wire   [3:0] MCInst2_MC2_v2_0;
  wire   [2:1] MCInst2_MC2_v1_3;
  wire   [3:0] MCInst2_MC2_v1_2;
  wire   [3:0] MCInst2_MC2_v1_1;
  wire   [3:0] MCInst2_MC2_v1_0;
  wire   [3:0] MCInst2_MC2_v0_3;
  wire   [3:0] MCInst2_MC2_v0_2;
  wire   [3:1] MCInst2_MC2_v0_1;
  wire   [3:1] MCInst2_MC2_v0_0;
  wire   [3:0] MCInst2_MC3_v3_3;
  wire   [3:0] MCInst2_MC3_v3_2;
  wire   [3:0] MCInst2_MC3_v3_1;
  wire   [2:1] MCInst2_MC3_v3_0;
  wire   [3:0] MCInst2_MC3_v2_3;
  wire   [3:0] MCInst2_MC3_v2_2;
  wire   [3:0] MCInst2_MC3_v2_1;
  wire   [3:0] MCInst2_MC3_v2_0;
  wire   [2:1] MCInst2_MC3_v1_3;
  wire   [3:0] MCInst2_MC3_v1_2;
  wire   [3:0] MCInst2_MC3_v1_1;
  wire   [3:0] MCInst2_MC3_v1_0;
  wire   [3:0] MCInst2_MC3_v0_3;
  wire   [3:0] MCInst2_MC3_v0_2;
  wire   [3:1] MCInst2_MC3_v0_1;
  wire   [3:1] MCInst2_MC3_v0_0;

  INV_X1 U4 ( .A(Error_0_), .ZN(ErrorFlag) );
  XOR2_X1 AddKeyXOR_XORInst_0_0_U1 ( .A(Plaintext[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR_XORInst_0_1_U1 ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR_XORInst_0_2_U1 ( .A(Plaintext[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR_XORInst_0_3_U1 ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR_XORInst_1_0_U1 ( .A(Plaintext[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR_XORInst_1_1_U1 ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR_XORInst_1_2_U1 ( .A(Plaintext[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR_XORInst_1_3_U1 ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR_XORInst_2_0_U1 ( .A(Plaintext[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR_XORInst_2_1_U1 ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR_XORInst_2_2_U1 ( .A(Plaintext[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR_XORInst_2_3_U1 ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR_XORInst_3_0_U1 ( .A(Plaintext[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR_XORInst_3_1_U1 ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR_XORInst_3_2_U1 ( .A(Plaintext[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR_XORInst_3_3_U1 ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR_XORInst_4_0_U1 ( .A(Plaintext[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR_XORInst_4_1_U1 ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR_XORInst_4_2_U1 ( .A(Plaintext[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR_XORInst_4_3_U1 ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR_XORInst_5_0_U1 ( .A(Plaintext[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR_XORInst_5_1_U1 ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR_XORInst_5_2_U1 ( .A(Plaintext[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR_XORInst_5_3_U1 ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR_XORInst_6_0_U1 ( .A(Plaintext[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR_XORInst_6_1_U1 ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR_XORInst_6_2_U1 ( .A(Plaintext[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR_XORInst_6_3_U1 ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR_XORInst_7_0_U1 ( .A(Plaintext[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR_XORInst_7_1_U1 ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR_XORInst_7_2_U1 ( .A(Plaintext[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR_XORInst_7_3_U1 ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR_XORInst_8_0_U1 ( .A(Plaintext[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR_XORInst_8_1_U1 ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR_XORInst_8_2_U1 ( .A(Plaintext[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR_XORInst_8_3_U1 ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR_XORInst_9_0_U1 ( .A(Plaintext[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR_XORInst_9_1_U1 ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR_XORInst_9_2_U1 ( .A(Plaintext[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR_XORInst_9_3_U1 ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  XOR2_X1 AddKeyXOR_XORInst_10_0_U1 ( .A(Plaintext[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X1 AddKeyXOR_XORInst_10_1_U1 ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X1 AddKeyXOR_XORInst_10_2_U1 ( .A(Plaintext[42]), .B(Key[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X1 AddKeyXOR_XORInst_10_3_U1 ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X1 AddKeyXOR_XORInst_11_0_U1 ( .A(Plaintext[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X1 AddKeyXOR_XORInst_11_1_U1 ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X1 AddKeyXOR_XORInst_11_2_U1 ( .A(Plaintext[46]), .B(Key[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X1 AddKeyXOR_XORInst_11_3_U1 ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X1 AddKeyXOR_XORInst_12_0_U1 ( .A(Plaintext[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR_XORInst_12_1_U1 ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR_XORInst_12_2_U1 ( .A(Plaintext[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR_XORInst_12_3_U1 ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR_XORInst_13_0_U1 ( .A(Plaintext[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR_XORInst_13_1_U1 ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR_XORInst_13_2_U1 ( .A(Plaintext[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR_XORInst_13_3_U1 ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR_XORInst_14_0_U1 ( .A(Plaintext[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR_XORInst_14_1_U1 ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR_XORInst_14_2_U1 ( .A(Plaintext[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR_XORInst_14_3_U1 ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR_XORInst_15_0_U1 ( .A(Plaintext[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR_XORInst_15_1_U1 ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR_XORInst_15_2_U1 ( .A(Plaintext[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR_XORInst_15_3_U1 ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_0_U4 ( .A1(AddRoundKeyOutput[2]), .A2(
        SubCellInst_LFInst_0_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U3 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_0_U2 ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .ZN(SubCellInst_LFInst_0_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_0_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_0_LFInst_0_n5), .B(SubCellInst_LFInst_0_LFInst_0_n7), .Z(MCInst_MC0_v3_2[3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n26), .A2(
        SubCellInst_LFInst_0_LFInst_1_n25), .ZN(MCInst_MC0_v3_0[2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n24), .A2(
        SubCellInst_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U8 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U7 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n21), .A2(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n20), .A2(
        SubCellInst_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n19), .A2(
        SubCellInst_LFInst_0_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U1 ( .A(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n25), .A2(
        SubCellInst_LFInst_0_LFInst_2_n28), .ZN(Red_MCInst_MC0_v3_1_0_) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U7 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_0_LFInst_2_n26), .B(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n22), .A2(
        SubCellInst_LFInst_0_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_2_U3 ( .A(AddRoundKeyOutput[2]), .B(
        SubCellInst_LFInst_0_LFInst_2_n23), .Z(
        SubCellInst_LFInst_0_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U9 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n23), .A2(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U7 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n23), .A2(
        SubCellInst_LFInst_0_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n20), .A2(
        SubCellInst_LFInst_0_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4 ( .A1(AddRoundKeyOutput[2]), .A2(
        AddRoundKeyOutput[0]), .ZN(SubCellInst_LFInst_0_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_0_LFInst_3_U3 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n26), .A2(
        SubCellInst_LFInst_0_LFInst_3_n25), .ZN(MCInst_MC0_v3_2[2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_0_U4 ( .A1(AddRoundKeyOutput[6]), .A2(
        SubCellInst_LFInst_1_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U3 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_0_U2 ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .ZN(SubCellInst_LFInst_1_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_1_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_1_LFInst_0_n5), .B(SubCellInst_LFInst_1_LFInst_0_n7), .Z(MCInst_MC3_v3_2[3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n26), .A2(
        SubCellInst_LFInst_1_LFInst_1_n25), .ZN(MCInst_MC3_v3_0[2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n24), .A2(
        SubCellInst_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U8 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U7 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n21), .A2(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n20), .A2(
        SubCellInst_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n19), .A2(
        SubCellInst_LFInst_1_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U2 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U1 ( .A(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n25), .A2(
        SubCellInst_LFInst_1_LFInst_2_n28), .ZN(Red_MCInst_MC3_v3_1_0_) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U7 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_1_LFInst_2_n26), .B(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n22), .A2(
        SubCellInst_LFInst_1_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_2_U3 ( .A(AddRoundKeyOutput[6]), .B(
        SubCellInst_LFInst_1_LFInst_2_n23), .Z(
        SubCellInst_LFInst_1_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U2 ( .A1(AddRoundKeyOutput[5]), .A2(
        AddRoundKeyOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U9 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n23), .A2(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U7 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n23), .A2(
        SubCellInst_LFInst_1_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n20), .A2(
        SubCellInst_LFInst_1_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4 ( .A1(AddRoundKeyOutput[6]), .A2(
        AddRoundKeyOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_1_LFInst_3_U3 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U2 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n26), .A2(
        SubCellInst_LFInst_1_LFInst_3_n25), .ZN(MCInst_MC3_v3_2[2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_0_U4 ( .A1(AddRoundKeyOutput[10]), .A2(
        SubCellInst_LFInst_2_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U3 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_0_U2 ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .ZN(SubCellInst_LFInst_2_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_2_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_2_LFInst_0_n5), .B(SubCellInst_LFInst_2_LFInst_0_n7), .Z(MCInst_MC2_v3_2[3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n26), .A2(
        SubCellInst_LFInst_2_LFInst_1_n25), .ZN(MCInst_MC2_v3_0[2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n24), .A2(
        SubCellInst_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U8 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U7 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n21), .A2(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n20), .A2(
        SubCellInst_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n19), .A2(
        SubCellInst_LFInst_2_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U2 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U1 ( .A(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n25), .A2(
        SubCellInst_LFInst_2_LFInst_2_n28), .ZN(Red_MCInst_MC2_v3_1_0_) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U7 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_2_LFInst_2_n26), .B(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n22), .A2(
        SubCellInst_LFInst_2_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_2_U3 ( .A(AddRoundKeyOutput[10]), .B(
        SubCellInst_LFInst_2_LFInst_2_n23), .Z(
        SubCellInst_LFInst_2_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U2 ( .A1(AddRoundKeyOutput[9]), .A2(
        AddRoundKeyOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U1 ( .A(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U9 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n23), .A2(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U7 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n23), .A2(
        SubCellInst_LFInst_2_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n20), .A2(
        SubCellInst_LFInst_2_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4 ( .A1(AddRoundKeyOutput[10]), .A2(
        AddRoundKeyOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_2_LFInst_3_U3 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U2 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n26), .A2(
        SubCellInst_LFInst_2_LFInst_3_n25), .ZN(MCInst_MC2_v3_2[2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_0_U4 ( .A1(AddRoundKeyOutput[14]), .A2(
        SubCellInst_LFInst_3_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U3 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_0_U2 ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .ZN(SubCellInst_LFInst_3_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_3_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_3_LFInst_0_n5), .B(SubCellInst_LFInst_3_LFInst_0_n7), .Z(MCInst_MC1_v3_2[3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n26), .A2(
        SubCellInst_LFInst_3_LFInst_1_n25), .ZN(MCInst_MC1_v3_0[2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n24), .A2(
        SubCellInst_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U8 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U7 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n21), .A2(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n20), .A2(
        SubCellInst_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n19), .A2(
        SubCellInst_LFInst_3_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U2 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U1 ( .A(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n25), .A2(
        SubCellInst_LFInst_3_LFInst_2_n28), .ZN(Red_MCInst_MC1_v3_1_0_) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U7 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_3_LFInst_2_n26), .B(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n22), .A2(
        SubCellInst_LFInst_3_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_2_U3 ( .A(AddRoundKeyOutput[14]), .B(
        SubCellInst_LFInst_3_LFInst_2_n23), .Z(
        SubCellInst_LFInst_3_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U2 ( .A1(AddRoundKeyOutput[13]), .A2(
        AddRoundKeyOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U1 ( .A(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U9 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n23), .A2(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U7 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n23), .A2(
        SubCellInst_LFInst_3_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n20), .A2(
        SubCellInst_LFInst_3_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4 ( .A1(AddRoundKeyOutput[14]), .A2(
        AddRoundKeyOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_3_LFInst_3_U3 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U2 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n26), .A2(
        SubCellInst_LFInst_3_LFInst_3_n25), .ZN(MCInst_MC1_v3_2[2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_0_U4 ( .A1(AddRoundKeyOutput[18]), .A2(
        SubCellInst_LFInst_4_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U3 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_0_U2 ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .ZN(SubCellInst_LFInst_4_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_4_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_4_LFInst_0_n5), .B(SubCellInst_LFInst_4_LFInst_0_n7), .Z(MCInst_MC1_v2_3[1]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n24), .A2(
        SubCellInst_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U9 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U8 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n21), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n20), .A2(
        SubCellInst_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U5 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n19), .A2(
        SubCellInst_LFInst_4_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U3 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U2 ( .A(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n26), .A2(
        SubCellInst_LFInst_4_LFInst_1_n25), .ZN(MCInst_MC1_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n25), .A2(
        SubCellInst_LFInst_4_LFInst_2_n28), .ZN(MCInst_MC1_v2_0[3]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U7 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_4_LFInst_2_n26), .B(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_2_U5 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n22), .A2(
        SubCellInst_LFInst_4_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_2_U3 ( .A(AddRoundKeyOutput[18]), .B(
        SubCellInst_LFInst_4_LFInst_2_n23), .Z(
        SubCellInst_LFInst_4_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U2 ( .A1(AddRoundKeyOutput[17]), .A2(
        AddRoundKeyOutput[16]), .ZN(SubCellInst_LFInst_4_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U1 ( .A(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U9 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n23), .A2(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_3_U7 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n23), .A2(
        SubCellInst_LFInst_4_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n20), .A2(
        SubCellInst_LFInst_4_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4 ( .A1(AddRoundKeyOutput[18]), .A2(
        AddRoundKeyOutput[16]), .ZN(SubCellInst_LFInst_4_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_4_LFInst_3_U3 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U2 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n26), .A2(
        SubCellInst_LFInst_4_LFInst_3_n25), .ZN(MCInst_MC1_v2_0[0]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_0_U4 ( .A1(AddRoundKeyOutput[22]), .A2(
        SubCellInst_LFInst_5_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U3 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_0_U2 ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .ZN(SubCellInst_LFInst_5_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_5_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_5_LFInst_0_n5), .B(SubCellInst_LFInst_5_LFInst_0_n7), .Z(MCInst_MC0_v2_3[1]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n24), .A2(
        SubCellInst_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U9 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U8 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n21), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n20), .A2(
        SubCellInst_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U5 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n19), .A2(
        SubCellInst_LFInst_5_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U3 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U2 ( .A(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n26), .A2(
        SubCellInst_LFInst_5_LFInst_1_n25), .ZN(MCInst_MC0_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n25), .A2(
        SubCellInst_LFInst_5_LFInst_2_n28), .ZN(MCInst_MC0_v2_0[3]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U7 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_5_LFInst_2_n26), .B(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_2_U5 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n22), .A2(
        SubCellInst_LFInst_5_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_2_U3 ( .A(AddRoundKeyOutput[22]), .B(
        SubCellInst_LFInst_5_LFInst_2_n23), .Z(
        SubCellInst_LFInst_5_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U2 ( .A1(AddRoundKeyOutput[21]), .A2(
        AddRoundKeyOutput[20]), .ZN(SubCellInst_LFInst_5_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U1 ( .A(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U9 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n23), .A2(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_3_U7 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n23), .A2(
        SubCellInst_LFInst_5_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n20), .A2(
        SubCellInst_LFInst_5_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4 ( .A1(AddRoundKeyOutput[22]), .A2(
        AddRoundKeyOutput[20]), .ZN(SubCellInst_LFInst_5_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_5_LFInst_3_U3 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U2 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n26), .A2(
        SubCellInst_LFInst_5_LFInst_3_n25), .ZN(MCInst_MC0_v2_0[0]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_0_U4 ( .A1(AddRoundKeyOutput[26]), .A2(
        SubCellInst_LFInst_6_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U3 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_0_U2 ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .ZN(SubCellInst_LFInst_6_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_6_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_6_LFInst_0_n5), .B(SubCellInst_LFInst_6_LFInst_0_n7), .Z(MCInst_MC3_v2_3[1]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n24), .A2(
        SubCellInst_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U9 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U8 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n21), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n20), .A2(
        SubCellInst_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U5 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n19), .A2(
        SubCellInst_LFInst_6_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U3 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U2 ( .A(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n26), .A2(
        SubCellInst_LFInst_6_LFInst_1_n25), .ZN(MCInst_MC3_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n25), .A2(
        SubCellInst_LFInst_6_LFInst_2_n28), .ZN(MCInst_MC3_v2_0[3]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U7 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_6_LFInst_2_n26), .B(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_2_U5 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n22), .A2(
        SubCellInst_LFInst_6_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_2_U3 ( .A(AddRoundKeyOutput[26]), .B(
        SubCellInst_LFInst_6_LFInst_2_n23), .Z(
        SubCellInst_LFInst_6_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U2 ( .A1(AddRoundKeyOutput[25]), .A2(
        AddRoundKeyOutput[24]), .ZN(SubCellInst_LFInst_6_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U1 ( .A(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U9 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n23), .A2(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_3_U7 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n23), .A2(
        SubCellInst_LFInst_6_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n20), .A2(
        SubCellInst_LFInst_6_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4 ( .A1(AddRoundKeyOutput[26]), .A2(
        AddRoundKeyOutput[24]), .ZN(SubCellInst_LFInst_6_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_6_LFInst_3_U3 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U2 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n26), .A2(
        SubCellInst_LFInst_6_LFInst_3_n25), .ZN(MCInst_MC3_v2_0[0]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_0_U4 ( .A1(AddRoundKeyOutput[30]), .A2(
        SubCellInst_LFInst_7_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U3 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_0_U2 ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .ZN(SubCellInst_LFInst_7_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_7_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_7_LFInst_0_n5), .B(SubCellInst_LFInst_7_LFInst_0_n7), .Z(MCInst_MC2_v2_3[1]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n24), .A2(
        SubCellInst_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U9 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U8 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n21), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n20), .A2(
        SubCellInst_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U5 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n19), .A2(
        SubCellInst_LFInst_7_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U3 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U2 ( .A(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n26), .A2(
        SubCellInst_LFInst_7_LFInst_1_n25), .ZN(MCInst_MC2_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n25), .A2(
        SubCellInst_LFInst_7_LFInst_2_n28), .ZN(MCInst_MC2_v2_0[3]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U7 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_7_LFInst_2_n26), .B(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_2_U5 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n22), .A2(
        SubCellInst_LFInst_7_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_2_U3 ( .A(AddRoundKeyOutput[30]), .B(
        SubCellInst_LFInst_7_LFInst_2_n23), .Z(
        SubCellInst_LFInst_7_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U2 ( .A1(AddRoundKeyOutput[29]), .A2(
        AddRoundKeyOutput[28]), .ZN(SubCellInst_LFInst_7_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U1 ( .A(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U9 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n23), .A2(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_3_U7 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n23), .A2(
        SubCellInst_LFInst_7_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n20), .A2(
        SubCellInst_LFInst_7_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4 ( .A1(AddRoundKeyOutput[30]), .A2(
        AddRoundKeyOutput[28]), .ZN(SubCellInst_LFInst_7_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_7_LFInst_3_U3 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U2 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n26), .A2(
        SubCellInst_LFInst_7_LFInst_3_n25), .ZN(MCInst_MC2_v2_0[0]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_0_U4 ( .A1(AddRoundKeyOutput[34]), .A2(
        SubCellInst_LFInst_8_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U3 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_0_U2 ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .ZN(SubCellInst_LFInst_8_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_8_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_8_LFInst_0_n5), .B(SubCellInst_LFInst_8_LFInst_0_n7), .Z(MCInst_MC2_v1_0[0]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n26), .A2(
        SubCellInst_LFInst_8_LFInst_1_n25), .ZN(MCInst_MC2_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n24), .A2(
        SubCellInst_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U8 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U7 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n21), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n20), .A2(
        SubCellInst_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n19), .A2(
        SubCellInst_LFInst_8_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U1 ( .A(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n25), .A2(
        SubCellInst_LFInst_8_LFInst_2_n28), .ZN(Red_MCInst_MC2_v1_1_0_) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U7 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_8_LFInst_2_n26), .B(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_2_U5 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n22), .A2(
        SubCellInst_LFInst_8_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U3 ( .A(AddRoundKeyOutput[34]), .B(
        SubCellInst_LFInst_8_LFInst_2_n23), .Z(
        SubCellInst_LFInst_8_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U2 ( .A1(AddRoundKeyOutput[33]), .A2(
        AddRoundKeyOutput[32]), .ZN(SubCellInst_LFInst_8_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U1 ( .A(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n26), .A2(
        SubCellInst_LFInst_8_LFInst_3_n25), .ZN(MCInst_MC2_v1_0[3]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U8 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n23), .A2(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U6 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n23), .A2(
        SubCellInst_LFInst_8_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n20), .A2(
        SubCellInst_LFInst_8_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U3 ( .A1(AddRoundKeyOutput[34]), .A2(
        AddRoundKeyOutput[32]), .ZN(SubCellInst_LFInst_8_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_8_LFInst_3_U2 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U1 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_0_U4 ( .A1(AddRoundKeyOutput[38]), .A2(
        SubCellInst_LFInst_9_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U3 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_0_U2 ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .ZN(SubCellInst_LFInst_9_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_9_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_9_LFInst_0_n5), .B(SubCellInst_LFInst_9_LFInst_0_n7), .Z(MCInst_MC1_v1_0[0]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n26), .A2(
        SubCellInst_LFInst_9_LFInst_1_n25), .ZN(MCInst_MC1_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n24), .A2(
        SubCellInst_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U8 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U7 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n21), .A2(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n20), .A2(
        SubCellInst_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n19), .A2(
        SubCellInst_LFInst_9_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U1 ( .A(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n25), .A2(
        SubCellInst_LFInst_9_LFInst_2_n28), .ZN(Red_MCInst_MC1_v1_1_0_) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U7 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_9_LFInst_2_n26), .B(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n22), .A2(
        SubCellInst_LFInst_9_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_2_U3 ( .A(AddRoundKeyOutput[38]), .B(
        SubCellInst_LFInst_9_LFInst_2_n23), .Z(
        SubCellInst_LFInst_9_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U2 ( .A1(AddRoundKeyOutput[37]), .A2(
        AddRoundKeyOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U1 ( .A(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n26), .A2(
        SubCellInst_LFInst_9_LFInst_3_n25), .ZN(MCInst_MC1_v1_0[3]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U8 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n23), .A2(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U6 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n23), .A2(
        SubCellInst_LFInst_9_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n20), .A2(
        SubCellInst_LFInst_9_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U3 ( .A1(AddRoundKeyOutput[38]), .A2(
        AddRoundKeyOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_9_LFInst_3_U2 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U1 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_0_U4 ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U3 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_0_U2 ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .ZN(SubCellInst_LFInst_10_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_10_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_10_LFInst_0_n5), .B(
        SubCellInst_LFInst_10_LFInst_0_n7), .Z(MCInst_MC0_v1_0[0]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n26), .A2(
        SubCellInst_LFInst_10_LFInst_1_n25), .ZN(MCInst_MC0_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n24), .A2(
        SubCellInst_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U8 ( .A1(AddRoundKeyOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U7 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n21), .A2(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n20), .A2(
        SubCellInst_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n19), .A2(
        SubCellInst_LFInst_10_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U1 ( .A(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n25), .A2(
        SubCellInst_LFInst_10_LFInst_2_n28), .ZN(Red_MCInst_MC0_v1_1_0_) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U7 ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_10_LFInst_2_n26), .B(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(AddRoundKeyOutput[40]), .A2(
        AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n22), .A2(
        SubCellInst_LFInst_10_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_2_U3 ( .A(AddRoundKeyOutput[42]), .B(
        SubCellInst_LFInst_10_LFInst_2_n23), .Z(
        SubCellInst_LFInst_10_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U2 ( .A1(AddRoundKeyOutput[41]), 
        .A2(AddRoundKeyOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U1 ( .A(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n26), .A2(
        SubCellInst_LFInst_10_LFInst_3_n25), .ZN(MCInst_MC0_v1_0[3]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U8 ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n23), .A2(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U6 ( .A1(AddRoundKeyOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n23), .A2(
        SubCellInst_LFInst_10_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n20), .A2(
        SubCellInst_LFInst_10_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U3 ( .A1(AddRoundKeyOutput[42]), .A2(
        AddRoundKeyOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_10_LFInst_3_U2 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U1 ( .A1(AddRoundKeyOutput[40]), .A2(
        AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_0_U4 ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U3 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_0_U2 ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .ZN(SubCellInst_LFInst_11_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_11_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_11_LFInst_0_n5), .B(
        SubCellInst_LFInst_11_LFInst_0_n7), .Z(MCInst_MC3_v1_0[0]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n26), .A2(
        SubCellInst_LFInst_11_LFInst_1_n25), .ZN(MCInst_MC3_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n24), .A2(
        SubCellInst_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U8 ( .A1(AddRoundKeyOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U7 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n21), .A2(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n20), .A2(
        SubCellInst_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n19), .A2(
        SubCellInst_LFInst_11_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U1 ( .A(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n25), .A2(
        SubCellInst_LFInst_11_LFInst_2_n28), .ZN(Red_MCInst_MC3_v1_1_0_) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U7 ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_11_LFInst_2_n26), .B(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(AddRoundKeyOutput[44]), .A2(
        AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n22), .A2(
        SubCellInst_LFInst_11_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_2_U3 ( .A(AddRoundKeyOutput[46]), .B(
        SubCellInst_LFInst_11_LFInst_2_n23), .Z(
        SubCellInst_LFInst_11_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U2 ( .A1(AddRoundKeyOutput[45]), 
        .A2(AddRoundKeyOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n26), .A2(
        SubCellInst_LFInst_11_LFInst_3_n25), .ZN(MCInst_MC3_v1_0[3]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U8 ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n23), .A2(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U6 ( .A1(AddRoundKeyOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n23), .A2(
        SubCellInst_LFInst_11_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n20), .A2(
        SubCellInst_LFInst_11_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U3 ( .A1(AddRoundKeyOutput[46]), .A2(
        AddRoundKeyOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_11_LFInst_3_U2 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U1 ( .A1(AddRoundKeyOutput[44]), .A2(
        AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_0_U4 ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U3 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_0_U2 ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .ZN(SubCellInst_LFInst_12_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_12_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_12_LFInst_0_n5), .B(
        SubCellInst_LFInst_12_LFInst_0_n7), .Z(Red_MCInst_MC3_v0_1_0_) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n26), .A2(
        SubCellInst_LFInst_12_LFInst_1_n25), .ZN(MCInst_MC3_v0_0[3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n24), .A2(
        SubCellInst_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U8 ( .A1(AddRoundKeyOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U7 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n21), .A2(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n20), .A2(
        SubCellInst_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n19), .A2(
        SubCellInst_LFInst_12_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U2 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U1 ( .A(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n25), .A2(
        SubCellInst_LFInst_12_LFInst_2_n28), .ZN(MCInst_MC3_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U7 ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_12_LFInst_2_n26), .B(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_2_U5 ( .A1(AddRoundKeyOutput[48]), .A2(
        AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n22), .A2(
        SubCellInst_LFInst_12_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U3 ( .A(AddRoundKeyOutput[50]), .B(
        SubCellInst_LFInst_12_LFInst_2_n23), .Z(
        SubCellInst_LFInst_12_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U2 ( .A1(AddRoundKeyOutput[49]), 
        .A2(AddRoundKeyOutput[48]), .ZN(SubCellInst_LFInst_12_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U1 ( .A(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U9 ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n23), .A2(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U7 ( .A1(AddRoundKeyOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n23), .A2(
        SubCellInst_LFInst_12_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n20), .A2(
        SubCellInst_LFInst_12_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U4 ( .A1(AddRoundKeyOutput[50]), .A2(
        AddRoundKeyOutput[48]), .ZN(SubCellInst_LFInst_12_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_12_LFInst_3_U3 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U2 ( .A1(AddRoundKeyOutput[48]), .A2(
        AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n26), .A2(
        SubCellInst_LFInst_12_LFInst_3_n25), .ZN(MCInst_MC3_v0_3[0]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_0_U4 ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U3 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_0_U2 ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .ZN(SubCellInst_LFInst_13_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_13_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_13_LFInst_0_n5), .B(
        SubCellInst_LFInst_13_LFInst_0_n7), .Z(Red_MCInst_MC2_v0_1_0_) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n26), .A2(
        SubCellInst_LFInst_13_LFInst_1_n25), .ZN(MCInst_MC2_v0_0[3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n24), .A2(
        SubCellInst_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U8 ( .A1(AddRoundKeyOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U7 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n21), .A2(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n20), .A2(
        SubCellInst_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n19), .A2(
        SubCellInst_LFInst_13_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U2 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U1 ( .A(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n25), .A2(
        SubCellInst_LFInst_13_LFInst_2_n28), .ZN(MCInst_MC2_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U7 ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_13_LFInst_2_n26), .B(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_2_U5 ( .A1(AddRoundKeyOutput[52]), .A2(
        AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n22), .A2(
        SubCellInst_LFInst_13_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_2_U3 ( .A(AddRoundKeyOutput[54]), .B(
        SubCellInst_LFInst_13_LFInst_2_n23), .Z(
        SubCellInst_LFInst_13_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U2 ( .A1(AddRoundKeyOutput[53]), 
        .A2(AddRoundKeyOutput[52]), .ZN(SubCellInst_LFInst_13_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U9 ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n23), .A2(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U7 ( .A1(AddRoundKeyOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n23), .A2(
        SubCellInst_LFInst_13_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n20), .A2(
        SubCellInst_LFInst_13_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U4 ( .A1(AddRoundKeyOutput[54]), .A2(
        AddRoundKeyOutput[52]), .ZN(SubCellInst_LFInst_13_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_13_LFInst_3_U3 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U2 ( .A1(AddRoundKeyOutput[52]), .A2(
        AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n26), .A2(
        SubCellInst_LFInst_13_LFInst_3_n25), .ZN(MCInst_MC2_v0_3[0]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_0_U4 ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U3 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_0_U2 ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .ZN(SubCellInst_LFInst_14_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_14_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_14_LFInst_0_n5), .B(
        SubCellInst_LFInst_14_LFInst_0_n7), .Z(Red_MCInst_MC1_v0_1_0_) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n26), .A2(
        SubCellInst_LFInst_14_LFInst_1_n25), .ZN(MCInst_MC1_v0_0[3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n24), .A2(
        SubCellInst_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U8 ( .A1(AddRoundKeyOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U7 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n21), .A2(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n20), .A2(
        SubCellInst_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n19), .A2(
        SubCellInst_LFInst_14_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U2 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U1 ( .A(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n25), .A2(
        SubCellInst_LFInst_14_LFInst_2_n28), .ZN(MCInst_MC1_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U7 ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_14_LFInst_2_n26), .B(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_2_U5 ( .A1(AddRoundKeyOutput[56]), .A2(
        AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n22), .A2(
        SubCellInst_LFInst_14_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U3 ( .A(AddRoundKeyOutput[58]), .B(
        SubCellInst_LFInst_14_LFInst_2_n23), .Z(
        SubCellInst_LFInst_14_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U2 ( .A1(AddRoundKeyOutput[57]), 
        .A2(AddRoundKeyOutput[56]), .ZN(SubCellInst_LFInst_14_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U1 ( .A(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U9 ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n23), .A2(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U7 ( .A1(AddRoundKeyOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n23), .A2(
        SubCellInst_LFInst_14_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n20), .A2(
        SubCellInst_LFInst_14_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U4 ( .A1(AddRoundKeyOutput[58]), .A2(
        AddRoundKeyOutput[56]), .ZN(SubCellInst_LFInst_14_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_14_LFInst_3_U3 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U2 ( .A1(AddRoundKeyOutput[56]), .A2(
        AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n26), .A2(
        SubCellInst_LFInst_14_LFInst_3_n25), .ZN(MCInst_MC1_v0_3[0]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_0_U4 ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U3 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n6) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_0_U2 ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .ZN(SubCellInst_LFInst_15_LFInst_0_n5) );
  XOR2_X2 SubCellInst_LFInst_15_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_15_LFInst_0_n5), .B(
        SubCellInst_LFInst_15_LFInst_0_n7), .Z(Red_MCInst_MC0_v0_1_0_) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n26), .A2(
        SubCellInst_LFInst_15_LFInst_1_n25), .ZN(MCInst_MC0_v0_0[3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n24), .A2(
        SubCellInst_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U8 ( .A1(AddRoundKeyOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U7 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n21), .A2(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n20), .A2(
        SubCellInst_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n19), .A2(
        SubCellInst_LFInst_15_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U2 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U1 ( .A(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n25), .A2(
        SubCellInst_LFInst_15_LFInst_2_n28), .ZN(MCInst_MC0_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U7 ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_15_LFInst_2_n26), .B(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_2_U5 ( .A1(AddRoundKeyOutput[60]), .A2(
        AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n22), .A2(
        SubCellInst_LFInst_15_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U3 ( .A(AddRoundKeyOutput[62]), .B(
        SubCellInst_LFInst_15_LFInst_2_n23), .Z(
        SubCellInst_LFInst_15_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U2 ( .A1(AddRoundKeyOutput[61]), 
        .A2(AddRoundKeyOutput[60]), .ZN(SubCellInst_LFInst_15_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U1 ( .A(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U9 ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n23), .A2(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U7 ( .A1(AddRoundKeyOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n23), .A2(
        SubCellInst_LFInst_15_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n20), .A2(
        SubCellInst_LFInst_15_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U4 ( .A1(AddRoundKeyOutput[62]), .A2(
        AddRoundKeyOutput[60]), .ZN(SubCellInst_LFInst_15_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_15_LFInst_3_U3 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U2 ( .A1(AddRoundKeyOutput[60]), .A2(
        AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n26), .A2(
        SubCellInst_LFInst_15_LFInst_3_n25), .ZN(MCInst_MC0_v0_3[0]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U2 ( .A(MCInst_MC0_v0_2Inst_0_n3), .B(
        MCInst_MC0_v0_3[0]), .ZN(MCInst_MC0_v0_2[0]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_0[3]), .ZN(MCInst_MC0_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v1_1Inst_0_U1 ( .A(Red_MCInst_MC0_v1_1_0_), .B(
        MCInst_MC0_v1_0[3]), .Z(MCInst_MC0_v1_1[0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U2 ( .A(MCInst_MC0_v1_2Inst_0_n3), .B(
        MCInst_MC0_v1_0[3]), .ZN(MCInst_MC0_v1_2[0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        Red_MCInst_MC0_v1_1_0_), .ZN(MCInst_MC0_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v2_1Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(MCInst_MC0_v2_1[0]) );
  XOR2_X1 MCInst_MC0_v2_2Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[0]), .Z(MCInst_MC0_v2_2[0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U3 ( .A(MCInst_MC0_v2_3Inst_0_n6), .B(
        MCInst_MC0_v2_3Inst_0_n5), .ZN(MCInst_MC0_v2_3[0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        MCInst_MC0_v2_0[0]), .ZN(MCInst_MC0_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC0_v2_3Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC0_v3_1Inst_0_U1 ( .A(Red_MCInst_MC0_v3_1_0_), .B(
        MCInst_MC0_v3_2[2]), .Z(MCInst_MC0_v3_1[0]) );
  XOR2_X1 MCInst_MC0_v3_2Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[2]), .Z(MCInst_MC0_v3_2[0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U2 ( .A(MCInst_MC0_v3_3Inst_0_n3), .B(
        MCInst_MC0_v3_2[2]), .ZN(MCInst_MC0_v3_3[0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[2]), .ZN(MCInst_MC0_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v0_0Inst_1_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v0_3[0]), .Z(MCInst_MC0_v0_0[1]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_1_U1 ( .A(MCInst_MC0_v0_0[3]), .B(
        MCInst_MC0_v0_3[3]), .Z(MCInst_MC0_v0_1[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U2 ( .A(MCInst_MC0_v0_2Inst_1_n3), .B(
        MCInst_MC0_v0_3[0]), .ZN(MCInst_MC0_v0_2[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_3[3]), .ZN(MCInst_MC0_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_3[0]), .Z(MCInst_MC0_v0_3[1]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_1_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        Red_MCInst_MC0_v1_1_0_), .Z(MCInst_MC0_v1_1[1]) );
  XOR2_X1 MCInst_MC0_v1_2Inst_1_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .Z(MCInst_MC0_v1_2[1]) );
  XOR2_X1 MCInst_MC0_v1_3Inst_1_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_0[3]), .Z(MCInst_MC0_v1_3[1]) );
  XOR2_X1 MCInst_MC0_v2_0Inst_1_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[0]), .Z(MCInst_MC0_v2_0[1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U2 ( .A(MCInst_MC0_v2_1Inst_1_n3), .B(
        MCInst_MC0_v2_0[0]), .ZN(MCInst_MC0_v2_1[1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U3 ( .A(MCInst_MC0_v2_2Inst_1_n6), .B(
        MCInst_MC0_v2_2Inst_1_n5), .ZN(MCInst_MC0_v2_2[1]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        MCInst_MC0_v2_0[0]), .ZN(MCInst_MC0_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC0_v2_2Inst_1_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC0_v3_0Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_2[2]), .Z(MCInst_MC0_v3_0[1]) );
  XOR2_X1 MCInst_MC0_v3_1Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_1_0_), .Z(MCInst_MC0_v3_1[1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U2 ( .A(MCInst_MC0_v3_3Inst_1_n3), .B(
        MCInst_MC0_v3_2[2]), .ZN(MCInst_MC0_v3_3[1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_1_0_), .ZN(MCInst_MC0_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_3[0]), .Z(MCInst_MC0_v0_0[2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_2_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v0_3[0]), .Z(MCInst_MC0_v0_1[2]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_2_U1 ( .A(MCInst_MC0_v0_0[3]), .B(
        MCInst_MC0_v0_3[0]), .Z(MCInst_MC0_v0_2[2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U2 ( .A(MCInst_MC0_v1_1Inst_2_n3), .B(
        MCInst_MC0_v1_0[3]), .ZN(MCInst_MC0_v1_1[2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U2 ( .A(MCInst_MC0_v1_2Inst_2_n3), .B(
        Red_MCInst_MC0_v1_1_0_), .ZN(MCInst_MC0_v1_2[2]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U2 ( .A(MCInst_MC0_v2_1Inst_2_n3), .B(
        MCInst_MC0_v2_0[0]), .ZN(MCInst_MC0_v2_1[2]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U2 ( .A(MCInst_MC0_v2_2Inst_2_n3), .B(
        MCInst_MC0_v2_0[0]), .ZN(MCInst_MC0_v2_2[2]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC0_v2_3Inst_2_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_3[2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U2 ( .A(MCInst_MC0_v3_1Inst_2_n3), .B(
        MCInst_MC0_v3_2[2]), .ZN(MCInst_MC0_v3_1[2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[2]), .ZN(MCInst_MC0_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC0_v3_3Inst_2_U1 ( .A(MCInst_MC0_v3_0[2]), .B(
        MCInst_MC0_v3_2[2]), .Z(MCInst_MC0_v3_3[2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_3_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_3[0]), .Z(MCInst_MC0_v0_1[3]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_3_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_3[3]), .Z(MCInst_MC0_v0_2[3]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_3_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        Red_MCInst_MC0_v1_1_0_), .Z(MCInst_MC0_v1_1[3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U3 ( .A(MCInst_MC0_v1_2Inst_3_n6), .B(
        MCInst_MC0_v1_2Inst_3_n5), .ZN(MCInst_MC0_v1_2[3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U2 ( .A(Red_MCInst_MC0_v1_1_0_), .B(
        MCInst_MC0_v1_0[3]), .ZN(MCInst_MC0_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC0_v1_2Inst_3_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .Z(MCInst_MC0_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC0_v2_1Inst_3_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[0]), .Z(MCInst_MC0_v2_1[3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U2 ( .A(MCInst_MC0_v2_2Inst_3_n3), .B(
        MCInst_MC0_v2_0[0]), .ZN(MCInst_MC0_v2_2[3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U2 ( .A(MCInst_MC0_v2_3Inst_3_n3), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_3[3]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .ZN(MCInst_MC0_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC0_v3_1Inst_3_U1 ( .A(MCInst_MC0_v3_0[2]), .B(
        Red_MCInst_MC0_v3_1_0_), .Z(MCInst_MC0_v3_1[3]) );
  XOR2_X1 MCInst_MC0_v3_3Inst_3_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_1_0_), .Z(MCInst_MC0_v3_3[3]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_0_n8), .B(MCInst_MC0_r0Inst_XORInst_0_0_n7), .ZN(MC_output[60]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_0[0]), .B(
        MCInst_MC0_v1_0[0]), .ZN(MCInst_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v3_2[2]), .Z(MCInst_MC0_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_1_n8), .B(MCInst_MC0_r0Inst_XORInst_0_1_n7), .ZN(MC_output[61]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_0[1]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_0[1]), .B(
        MCInst_MC0_v3_0[1]), .Z(MCInst_MC0_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_2_n8), .B(MCInst_MC0_r0Inst_XORInst_0_2_n7), .ZN(MC_output[62]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_0[2]), .B(
        Red_MCInst_MC0_v1_1_0_), .ZN(MCInst_MC0_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_0[2]), .B(
        MCInst_MC0_v3_0[2]), .Z(MCInst_MC0_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_3_n8), .B(MCInst_MC0_r0Inst_XORInst_0_3_n7), .ZN(MC_output[63]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        MCInst_MC0_v1_0[3]), .ZN(MCInst_MC0_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_0[3]), .B(
        Red_MCInst_MC0_v3_1_0_), .Z(MCInst_MC0_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_0_n8), .B(MCInst_MC0_r1Inst_XORInst_0_0_n7), .ZN(MC_output[44]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_1[0]), .B(
        MCInst_MC0_v1_1[0]), .ZN(MCInst_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_0[3]), .B(
        MCInst_MC0_v3_1[0]), .Z(MCInst_MC0_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_1_n8), .B(MCInst_MC0_r1Inst_XORInst_0_1_n7), .ZN(MC_output[45]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v1_1[1]), .ZN(MCInst_MC0_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_1[1]), .B(
        MCInst_MC0_v3_1[1]), .Z(MCInst_MC0_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_2_n8), .B(MCInst_MC0_r1Inst_XORInst_0_2_n7), .ZN(MC_output[46]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_1[2]), .B(
        MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_1[2]), .B(
        MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_3_n8), .B(MCInst_MC0_r1Inst_XORInst_0_3_n7), .ZN(MC_output[47]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_1[3]), .B(
        MCInst_MC0_v1_1[3]), .ZN(MCInst_MC0_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_1[3]), .B(
        MCInst_MC0_v3_1[3]), .Z(MCInst_MC0_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_0_n8), .B(MCInst_MC0_r2Inst_XORInst_0_0_n7), .ZN(MC_output[28]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_2[0]), .B(
        MCInst_MC0_v1_2[0]), .ZN(MCInst_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_2[0]), .B(
        MCInst_MC0_v3_2[0]), .Z(MCInst_MC0_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_1_n8), .B(MCInst_MC0_r2Inst_XORInst_0_1_n7), .ZN(MC_output[29]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_2[1]), .B(
        MCInst_MC0_v1_2[1]), .ZN(MCInst_MC0_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_2[1]), .B(
        Red_MCInst_MC0_v3_1_0_), .Z(MCInst_MC0_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_2_n8), .B(MCInst_MC0_r2Inst_XORInst_0_2_n7), .ZN(MC_output[30]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_2[2]), .B(
        MCInst_MC0_v1_2[2]), .ZN(MCInst_MC0_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_2[2]), .Z(MCInst_MC0_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_3_n8), .B(MCInst_MC0_r2Inst_XORInst_0_3_n7), .ZN(MC_output[31]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_2[3]), .B(
        MCInst_MC0_v1_2[3]), .ZN(MCInst_MC0_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_2[3]), .B(
        MCInst_MC0_v3_2[3]), .Z(MCInst_MC0_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_0_n8), .B(MCInst_MC0_r3Inst_XORInst_0_0_n7), .ZN(MC_output[12]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_3[0]), .B(
        MCInst_MC0_v1_0[3]), .ZN(MCInst_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_3[0]), .B(
        MCInst_MC0_v3_3[0]), .Z(MCInst_MC0_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_1_n8), .B(MCInst_MC0_r3Inst_XORInst_0_1_n7), .ZN(MC_output[13]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v1_3[1]), .ZN(MCInst_MC0_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_3[1]), .B(
        MCInst_MC0_v3_3[1]), .Z(MCInst_MC0_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_2_n8), .B(MCInst_MC0_r3Inst_XORInst_0_2_n7), .ZN(MC_output[14]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_3[2]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_0[3]), .B(
        MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_3_n8), .B(MCInst_MC0_r3Inst_XORInst_0_3_n7), .ZN(MC_output[15]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_3[3]), .B(
        Red_MCInst_MC0_v1_1_0_), .ZN(MCInst_MC0_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v3_3[3]), .Z(MCInst_MC0_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U2 ( .A(MCInst_MC1_v0_2Inst_0_n3), .B(
        MCInst_MC1_v0_3[0]), .ZN(MCInst_MC1_v0_2[0]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_0[3]), .ZN(MCInst_MC1_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v1_1Inst_0_U1 ( .A(Red_MCInst_MC1_v1_1_0_), .B(
        MCInst_MC1_v1_0[3]), .Z(MCInst_MC1_v1_1[0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U2 ( .A(MCInst_MC1_v1_2Inst_0_n3), .B(
        MCInst_MC1_v1_0[3]), .ZN(MCInst_MC1_v1_2[0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        Red_MCInst_MC1_v1_1_0_), .ZN(MCInst_MC1_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v2_1Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(MCInst_MC1_v2_1[0]) );
  XOR2_X1 MCInst_MC1_v2_2Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[0]), .Z(MCInst_MC1_v2_2[0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U3 ( .A(MCInst_MC1_v2_3Inst_0_n6), .B(
        MCInst_MC1_v2_3Inst_0_n5), .ZN(MCInst_MC1_v2_3[0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        MCInst_MC1_v2_0[0]), .ZN(MCInst_MC1_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC1_v2_3Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC1_v3_1Inst_0_U1 ( .A(Red_MCInst_MC1_v3_1_0_), .B(
        MCInst_MC1_v3_2[2]), .Z(MCInst_MC1_v3_1[0]) );
  XOR2_X1 MCInst_MC1_v3_2Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[2]), .Z(MCInst_MC1_v3_2[0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U2 ( .A(MCInst_MC1_v3_3Inst_0_n3), .B(
        MCInst_MC1_v3_2[2]), .ZN(MCInst_MC1_v3_3[0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[2]), .ZN(MCInst_MC1_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v0_0Inst_1_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v0_3[0]), .Z(MCInst_MC1_v0_0[1]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_1_U1 ( .A(MCInst_MC1_v0_0[3]), .B(
        MCInst_MC1_v0_3[3]), .Z(MCInst_MC1_v0_1[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U2 ( .A(MCInst_MC1_v0_2Inst_1_n3), .B(
        MCInst_MC1_v0_3[0]), .ZN(MCInst_MC1_v0_2[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_3[3]), .ZN(MCInst_MC1_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_3[0]), .Z(MCInst_MC1_v0_3[1]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_1_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        Red_MCInst_MC1_v1_1_0_), .Z(MCInst_MC1_v1_1[1]) );
  XOR2_X1 MCInst_MC1_v1_2Inst_1_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .Z(MCInst_MC1_v1_2[1]) );
  XOR2_X1 MCInst_MC1_v1_3Inst_1_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_0[3]), .Z(MCInst_MC1_v1_3[1]) );
  XOR2_X1 MCInst_MC1_v2_0Inst_1_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[0]), .Z(MCInst_MC1_v2_0[1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U2 ( .A(MCInst_MC1_v2_1Inst_1_n3), .B(
        MCInst_MC1_v2_0[0]), .ZN(MCInst_MC1_v2_1[1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U3 ( .A(MCInst_MC1_v2_2Inst_1_n6), .B(
        MCInst_MC1_v2_2Inst_1_n5), .ZN(MCInst_MC1_v2_2[1]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        MCInst_MC1_v2_0[0]), .ZN(MCInst_MC1_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC1_v2_2Inst_1_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC1_v3_0Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_2[2]), .Z(MCInst_MC1_v3_0[1]) );
  XOR2_X1 MCInst_MC1_v3_1Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_1_0_), .Z(MCInst_MC1_v3_1[1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U2 ( .A(MCInst_MC1_v3_3Inst_1_n3), .B(
        MCInst_MC1_v3_2[2]), .ZN(MCInst_MC1_v3_3[1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_1_0_), .ZN(MCInst_MC1_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_3[0]), .Z(MCInst_MC1_v0_0[2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_2_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v0_3[0]), .Z(MCInst_MC1_v0_1[2]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_2_U1 ( .A(MCInst_MC1_v0_0[3]), .B(
        MCInst_MC1_v0_3[0]), .Z(MCInst_MC1_v0_2[2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U2 ( .A(MCInst_MC1_v1_1Inst_2_n3), .B(
        MCInst_MC1_v1_0[3]), .ZN(MCInst_MC1_v1_1[2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U2 ( .A(MCInst_MC1_v1_2Inst_2_n3), .B(
        Red_MCInst_MC1_v1_1_0_), .ZN(MCInst_MC1_v1_2[2]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U2 ( .A(MCInst_MC1_v2_1Inst_2_n3), .B(
        MCInst_MC1_v2_0[0]), .ZN(MCInst_MC1_v2_1[2]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U2 ( .A(MCInst_MC1_v2_2Inst_2_n3), .B(
        MCInst_MC1_v2_0[0]), .ZN(MCInst_MC1_v2_2[2]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC1_v2_3Inst_2_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_3[2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U2 ( .A(MCInst_MC1_v3_1Inst_2_n3), .B(
        MCInst_MC1_v3_2[2]), .ZN(MCInst_MC1_v3_1[2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[2]), .ZN(MCInst_MC1_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC1_v3_3Inst_2_U1 ( .A(MCInst_MC1_v3_0[2]), .B(
        MCInst_MC1_v3_2[2]), .Z(MCInst_MC1_v3_3[2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_3_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_3[0]), .Z(MCInst_MC1_v0_1[3]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_3_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_3[3]), .Z(MCInst_MC1_v0_2[3]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_3_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        Red_MCInst_MC1_v1_1_0_), .Z(MCInst_MC1_v1_1[3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U3 ( .A(MCInst_MC1_v1_2Inst_3_n6), .B(
        MCInst_MC1_v1_2Inst_3_n5), .ZN(MCInst_MC1_v1_2[3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U2 ( .A(Red_MCInst_MC1_v1_1_0_), .B(
        MCInst_MC1_v1_0[3]), .ZN(MCInst_MC1_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC1_v1_2Inst_3_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .Z(MCInst_MC1_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC1_v2_1Inst_3_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[0]), .Z(MCInst_MC1_v2_1[3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U2 ( .A(MCInst_MC1_v2_2Inst_3_n3), .B(
        MCInst_MC1_v2_0[0]), .ZN(MCInst_MC1_v2_2[3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U2 ( .A(MCInst_MC1_v2_3Inst_3_n3), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_3[3]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .ZN(MCInst_MC1_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC1_v3_1Inst_3_U1 ( .A(MCInst_MC1_v3_0[2]), .B(
        Red_MCInst_MC1_v3_1_0_), .Z(MCInst_MC1_v3_1[3]) );
  XOR2_X1 MCInst_MC1_v3_3Inst_3_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_1_0_), .Z(MCInst_MC1_v3_3[3]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_0_n8), .B(MCInst_MC1_r0Inst_XORInst_0_0_n7), .ZN(MC_output[56]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_0[0]), .B(
        MCInst_MC1_v1_0[0]), .ZN(MCInst_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v3_2[2]), .Z(MCInst_MC1_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_1_n8), .B(MCInst_MC1_r0Inst_XORInst_0_1_n7), .ZN(MC_output[57]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_0[1]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_0[1]), .B(
        MCInst_MC1_v3_0[1]), .Z(MCInst_MC1_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_2_n8), .B(MCInst_MC1_r0Inst_XORInst_0_2_n7), .ZN(MC_output[58]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_0[2]), .B(
        Red_MCInst_MC1_v1_1_0_), .ZN(MCInst_MC1_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_0[2]), .B(
        MCInst_MC1_v3_0[2]), .Z(MCInst_MC1_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_3_n8), .B(MCInst_MC1_r0Inst_XORInst_0_3_n7), .ZN(MC_output[59]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        MCInst_MC1_v1_0[3]), .ZN(MCInst_MC1_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_0[3]), .B(
        Red_MCInst_MC1_v3_1_0_), .Z(MCInst_MC1_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_0_n8), .B(MCInst_MC1_r1Inst_XORInst_0_0_n7), .ZN(MC_output[40]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_1[0]), .B(
        MCInst_MC1_v1_1[0]), .ZN(MCInst_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_0[3]), .B(
        MCInst_MC1_v3_1[0]), .Z(MCInst_MC1_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_1_n8), .B(MCInst_MC1_r1Inst_XORInst_0_1_n7), .ZN(MC_output[41]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v1_1[1]), .ZN(MCInst_MC1_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_1[1]), .B(
        MCInst_MC1_v3_1[1]), .Z(MCInst_MC1_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_2_n8), .B(MCInst_MC1_r1Inst_XORInst_0_2_n7), .ZN(MC_output[42]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_1[2]), .B(
        MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_1[2]), .B(
        MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_3_n8), .B(MCInst_MC1_r1Inst_XORInst_0_3_n7), .ZN(MC_output[43]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_1[3]), .B(
        MCInst_MC1_v1_1[3]), .ZN(MCInst_MC1_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_1[3]), .B(
        MCInst_MC1_v3_1[3]), .Z(MCInst_MC1_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_0_n8), .B(MCInst_MC1_r2Inst_XORInst_0_0_n7), .ZN(MC_output[24]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_2[0]), .B(
        MCInst_MC1_v1_2[0]), .ZN(MCInst_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_2[0]), .B(
        MCInst_MC1_v3_2[0]), .Z(MCInst_MC1_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_1_n8), .B(MCInst_MC1_r2Inst_XORInst_0_1_n7), .ZN(MC_output[25]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_2[1]), .B(
        MCInst_MC1_v1_2[1]), .ZN(MCInst_MC1_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_2[1]), .B(
        Red_MCInst_MC1_v3_1_0_), .Z(MCInst_MC1_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_2_n8), .B(MCInst_MC1_r2Inst_XORInst_0_2_n7), .ZN(MC_output[26]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_2[2]), .B(
        MCInst_MC1_v1_2[2]), .ZN(MCInst_MC1_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_2[2]), .Z(MCInst_MC1_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_3_n8), .B(MCInst_MC1_r2Inst_XORInst_0_3_n7), .ZN(MC_output[27]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_2[3]), .B(
        MCInst_MC1_v1_2[3]), .ZN(MCInst_MC1_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_2[3]), .B(
        MCInst_MC1_v3_2[3]), .Z(MCInst_MC1_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_0_n8), .B(MCInst_MC1_r3Inst_XORInst_0_0_n7), .ZN(MC_output[8]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_3[0]), .B(
        MCInst_MC1_v1_0[3]), .ZN(MCInst_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_3[0]), .B(
        MCInst_MC1_v3_3[0]), .Z(MCInst_MC1_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_1_n8), .B(MCInst_MC1_r3Inst_XORInst_0_1_n7), .ZN(MC_output[9]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v1_3[1]), .ZN(MCInst_MC1_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_3[1]), .B(
        MCInst_MC1_v3_3[1]), .Z(MCInst_MC1_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_2_n8), .B(MCInst_MC1_r3Inst_XORInst_0_2_n7), .ZN(MC_output[10]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_3[2]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_0[3]), .B(
        MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_3_n8), .B(MCInst_MC1_r3Inst_XORInst_0_3_n7), .ZN(MC_output[11]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_3[3]), .B(
        Red_MCInst_MC1_v1_1_0_), .ZN(MCInst_MC1_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v3_3[3]), .Z(MCInst_MC1_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U2 ( .A(MCInst_MC2_v0_2Inst_0_n3), .B(
        MCInst_MC2_v0_3[0]), .ZN(MCInst_MC2_v0_2[0]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_0[3]), .ZN(MCInst_MC2_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v1_1Inst_0_U1 ( .A(Red_MCInst_MC2_v1_1_0_), .B(
        MCInst_MC2_v1_0[3]), .Z(MCInst_MC2_v1_1[0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U2 ( .A(MCInst_MC2_v1_2Inst_0_n3), .B(
        MCInst_MC2_v1_0[3]), .ZN(MCInst_MC2_v1_2[0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        Red_MCInst_MC2_v1_1_0_), .ZN(MCInst_MC2_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v2_1Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(MCInst_MC2_v2_1[0]) );
  XOR2_X1 MCInst_MC2_v2_2Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[0]), .Z(MCInst_MC2_v2_2[0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U3 ( .A(MCInst_MC2_v2_3Inst_0_n6), .B(
        MCInst_MC2_v2_3Inst_0_n5), .ZN(MCInst_MC2_v2_3[0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        MCInst_MC2_v2_0[0]), .ZN(MCInst_MC2_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC2_v2_3Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC2_v3_1Inst_0_U1 ( .A(Red_MCInst_MC2_v3_1_0_), .B(
        MCInst_MC2_v3_2[2]), .Z(MCInst_MC2_v3_1[0]) );
  XOR2_X1 MCInst_MC2_v3_2Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[2]), .Z(MCInst_MC2_v3_2[0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U2 ( .A(MCInst_MC2_v3_3Inst_0_n3), .B(
        MCInst_MC2_v3_2[2]), .ZN(MCInst_MC2_v3_3[0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[2]), .ZN(MCInst_MC2_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v0_0Inst_1_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v0_3[0]), .Z(MCInst_MC2_v0_0[1]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_1_U1 ( .A(MCInst_MC2_v0_0[3]), .B(
        MCInst_MC2_v0_3[3]), .Z(MCInst_MC2_v0_1[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U2 ( .A(MCInst_MC2_v0_2Inst_1_n3), .B(
        MCInst_MC2_v0_3[0]), .ZN(MCInst_MC2_v0_2[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_3[3]), .ZN(MCInst_MC2_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_3[0]), .Z(MCInst_MC2_v0_3[1]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_1_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        Red_MCInst_MC2_v1_1_0_), .Z(MCInst_MC2_v1_1[1]) );
  XOR2_X1 MCInst_MC2_v1_2Inst_1_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .Z(MCInst_MC2_v1_2[1]) );
  XOR2_X1 MCInst_MC2_v1_3Inst_1_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_0[3]), .Z(MCInst_MC2_v1_3[1]) );
  XOR2_X1 MCInst_MC2_v2_0Inst_1_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[0]), .Z(MCInst_MC2_v2_0[1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U2 ( .A(MCInst_MC2_v2_1Inst_1_n3), .B(
        MCInst_MC2_v2_0[0]), .ZN(MCInst_MC2_v2_1[1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U3 ( .A(MCInst_MC2_v2_2Inst_1_n6), .B(
        MCInst_MC2_v2_2Inst_1_n5), .ZN(MCInst_MC2_v2_2[1]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        MCInst_MC2_v2_0[0]), .ZN(MCInst_MC2_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC2_v2_2Inst_1_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC2_v3_0Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_2[2]), .Z(MCInst_MC2_v3_0[1]) );
  XOR2_X1 MCInst_MC2_v3_1Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_1_0_), .Z(MCInst_MC2_v3_1[1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U2 ( .A(MCInst_MC2_v3_3Inst_1_n3), .B(
        MCInst_MC2_v3_2[2]), .ZN(MCInst_MC2_v3_3[1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_1_0_), .ZN(MCInst_MC2_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_3[0]), .Z(MCInst_MC2_v0_0[2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_2_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v0_3[0]), .Z(MCInst_MC2_v0_1[2]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_2_U1 ( .A(MCInst_MC2_v0_0[3]), .B(
        MCInst_MC2_v0_3[0]), .Z(MCInst_MC2_v0_2[2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U2 ( .A(MCInst_MC2_v1_1Inst_2_n3), .B(
        MCInst_MC2_v1_0[3]), .ZN(MCInst_MC2_v1_1[2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U2 ( .A(MCInst_MC2_v1_2Inst_2_n3), .B(
        Red_MCInst_MC2_v1_1_0_), .ZN(MCInst_MC2_v1_2[2]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U2 ( .A(MCInst_MC2_v2_1Inst_2_n3), .B(
        MCInst_MC2_v2_0[0]), .ZN(MCInst_MC2_v2_1[2]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U2 ( .A(MCInst_MC2_v2_2Inst_2_n3), .B(
        MCInst_MC2_v2_0[0]), .ZN(MCInst_MC2_v2_2[2]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC2_v2_3Inst_2_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_3[2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U2 ( .A(MCInst_MC2_v3_1Inst_2_n3), .B(
        MCInst_MC2_v3_2[2]), .ZN(MCInst_MC2_v3_1[2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[2]), .ZN(MCInst_MC2_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC2_v3_3Inst_2_U1 ( .A(MCInst_MC2_v3_0[2]), .B(
        MCInst_MC2_v3_2[2]), .Z(MCInst_MC2_v3_3[2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_3_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_3[0]), .Z(MCInst_MC2_v0_1[3]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_3_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_3[3]), .Z(MCInst_MC2_v0_2[3]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_3_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        Red_MCInst_MC2_v1_1_0_), .Z(MCInst_MC2_v1_1[3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U3 ( .A(MCInst_MC2_v1_2Inst_3_n6), .B(
        MCInst_MC2_v1_2Inst_3_n5), .ZN(MCInst_MC2_v1_2[3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U2 ( .A(Red_MCInst_MC2_v1_1_0_), .B(
        MCInst_MC2_v1_0[3]), .ZN(MCInst_MC2_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC2_v1_2Inst_3_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .Z(MCInst_MC2_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC2_v2_1Inst_3_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[0]), .Z(MCInst_MC2_v2_1[3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U2 ( .A(MCInst_MC2_v2_2Inst_3_n3), .B(
        MCInst_MC2_v2_0[0]), .ZN(MCInst_MC2_v2_2[3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U2 ( .A(MCInst_MC2_v2_3Inst_3_n3), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_3[3]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .ZN(MCInst_MC2_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC2_v3_1Inst_3_U1 ( .A(MCInst_MC2_v3_0[2]), .B(
        Red_MCInst_MC2_v3_1_0_), .Z(MCInst_MC2_v3_1[3]) );
  XOR2_X1 MCInst_MC2_v3_3Inst_3_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_1_0_), .Z(MCInst_MC2_v3_3[3]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_0_n8), .B(MCInst_MC2_r0Inst_XORInst_0_0_n7), .ZN(MC_output[52]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_0[0]), .B(
        MCInst_MC2_v1_0[0]), .ZN(MCInst_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v3_2[2]), .Z(MCInst_MC2_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_1_n8), .B(MCInst_MC2_r0Inst_XORInst_0_1_n7), .ZN(MC_output[53]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_0[1]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_0[1]), .B(
        MCInst_MC2_v3_0[1]), .Z(MCInst_MC2_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_2_n8), .B(MCInst_MC2_r0Inst_XORInst_0_2_n7), .ZN(MC_output[54]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_0[2]), .B(
        Red_MCInst_MC2_v1_1_0_), .ZN(MCInst_MC2_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_0[2]), .B(
        MCInst_MC2_v3_0[2]), .Z(MCInst_MC2_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_3_n8), .B(MCInst_MC2_r0Inst_XORInst_0_3_n7), .ZN(MC_output[55]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        MCInst_MC2_v1_0[3]), .ZN(MCInst_MC2_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_0[3]), .B(
        Red_MCInst_MC2_v3_1_0_), .Z(MCInst_MC2_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_0_n8), .B(MCInst_MC2_r1Inst_XORInst_0_0_n7), .ZN(MC_output[36]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_1[0]), .B(
        MCInst_MC2_v1_1[0]), .ZN(MCInst_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_0[3]), .B(
        MCInst_MC2_v3_1[0]), .Z(MCInst_MC2_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_1_n8), .B(MCInst_MC2_r1Inst_XORInst_0_1_n7), .ZN(MC_output[37]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v1_1[1]), .ZN(MCInst_MC2_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_1[1]), .B(
        MCInst_MC2_v3_1[1]), .Z(MCInst_MC2_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_2_n8), .B(MCInst_MC2_r1Inst_XORInst_0_2_n7), .ZN(MC_output[38]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_1[2]), .B(
        MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_1[2]), .B(
        MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_3_n8), .B(MCInst_MC2_r1Inst_XORInst_0_3_n7), .ZN(MC_output[39]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_1[3]), .B(
        MCInst_MC2_v1_1[3]), .ZN(MCInst_MC2_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_1[3]), .B(
        MCInst_MC2_v3_1[3]), .Z(MCInst_MC2_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_0_n8), .B(MCInst_MC2_r2Inst_XORInst_0_0_n7), .ZN(MC_output[20]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_2[0]), .B(
        MCInst_MC2_v1_2[0]), .ZN(MCInst_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_2[0]), .B(
        MCInst_MC2_v3_2[0]), .Z(MCInst_MC2_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_1_n8), .B(MCInst_MC2_r2Inst_XORInst_0_1_n7), .ZN(MC_output[21]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_2[1]), .B(
        MCInst_MC2_v1_2[1]), .ZN(MCInst_MC2_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_2[1]), .B(
        Red_MCInst_MC2_v3_1_0_), .Z(MCInst_MC2_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_2_n8), .B(MCInst_MC2_r2Inst_XORInst_0_2_n7), .ZN(MC_output[22]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_2[2]), .B(
        MCInst_MC2_v1_2[2]), .ZN(MCInst_MC2_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_2[2]), .Z(MCInst_MC2_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_3_n8), .B(MCInst_MC2_r2Inst_XORInst_0_3_n7), .ZN(MC_output[23]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_2[3]), .B(
        MCInst_MC2_v1_2[3]), .ZN(MCInst_MC2_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_2[3]), .B(
        MCInst_MC2_v3_2[3]), .Z(MCInst_MC2_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_0_n8), .B(MCInst_MC2_r3Inst_XORInst_0_0_n7), .ZN(MC_output[4]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_3[0]), .B(
        MCInst_MC2_v1_0[3]), .ZN(MCInst_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_3[0]), .B(
        MCInst_MC2_v3_3[0]), .Z(MCInst_MC2_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_1_n8), .B(MCInst_MC2_r3Inst_XORInst_0_1_n7), .ZN(MC_output[5]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v1_3[1]), .ZN(MCInst_MC2_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_3[1]), .B(
        MCInst_MC2_v3_3[1]), .Z(MCInst_MC2_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_2_n8), .B(MCInst_MC2_r3Inst_XORInst_0_2_n7), .ZN(MC_output[6]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_3[2]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_0[3]), .B(
        MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_3_n8), .B(MCInst_MC2_r3Inst_XORInst_0_3_n7), .ZN(MC_output[7]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_3[3]), .B(
        Red_MCInst_MC2_v1_1_0_), .ZN(MCInst_MC2_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v3_3[3]), .Z(MCInst_MC2_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U2 ( .A(MCInst_MC3_v0_2Inst_0_n3), .B(
        MCInst_MC3_v0_3[0]), .ZN(MCInst_MC3_v0_2[0]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_0[3]), .ZN(MCInst_MC3_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v1_1Inst_0_U1 ( .A(Red_MCInst_MC3_v1_1_0_), .B(
        MCInst_MC3_v1_0[3]), .Z(MCInst_MC3_v1_1[0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U2 ( .A(MCInst_MC3_v1_2Inst_0_n3), .B(
        MCInst_MC3_v1_0[3]), .ZN(MCInst_MC3_v1_2[0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        Red_MCInst_MC3_v1_1_0_), .ZN(MCInst_MC3_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v2_1Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(MCInst_MC3_v2_1[0]) );
  XOR2_X1 MCInst_MC3_v2_2Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[0]), .Z(MCInst_MC3_v2_2[0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U3 ( .A(MCInst_MC3_v2_3Inst_0_n6), .B(
        MCInst_MC3_v2_3Inst_0_n5), .ZN(MCInst_MC3_v2_3[0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        MCInst_MC3_v2_0[0]), .ZN(MCInst_MC3_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC3_v2_3Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC3_v3_1Inst_0_U1 ( .A(Red_MCInst_MC3_v3_1_0_), .B(
        MCInst_MC3_v3_2[2]), .Z(MCInst_MC3_v3_1[0]) );
  XOR2_X1 MCInst_MC3_v3_2Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[2]), .Z(MCInst_MC3_v3_2[0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U2 ( .A(MCInst_MC3_v3_3Inst_0_n3), .B(
        MCInst_MC3_v3_2[2]), .ZN(MCInst_MC3_v3_3[0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[2]), .ZN(MCInst_MC3_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v0_0Inst_1_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v0_3[0]), .Z(MCInst_MC3_v0_0[1]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_1_U1 ( .A(MCInst_MC3_v0_0[3]), .B(
        MCInst_MC3_v0_3[3]), .Z(MCInst_MC3_v0_1[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U2 ( .A(MCInst_MC3_v0_2Inst_1_n3), .B(
        MCInst_MC3_v0_3[0]), .ZN(MCInst_MC3_v0_2[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_3[3]), .ZN(MCInst_MC3_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_3[0]), .Z(MCInst_MC3_v0_3[1]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_1_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        Red_MCInst_MC3_v1_1_0_), .Z(MCInst_MC3_v1_1[1]) );
  XOR2_X1 MCInst_MC3_v1_2Inst_1_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .Z(MCInst_MC3_v1_2[1]) );
  XOR2_X1 MCInst_MC3_v1_3Inst_1_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_0[3]), .Z(MCInst_MC3_v1_3[1]) );
  XOR2_X1 MCInst_MC3_v2_0Inst_1_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[0]), .Z(MCInst_MC3_v2_0[1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U2 ( .A(MCInst_MC3_v2_1Inst_1_n3), .B(
        MCInst_MC3_v2_0[0]), .ZN(MCInst_MC3_v2_1[1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U3 ( .A(MCInst_MC3_v2_2Inst_1_n6), .B(
        MCInst_MC3_v2_2Inst_1_n5), .ZN(MCInst_MC3_v2_2[1]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        MCInst_MC3_v2_0[0]), .ZN(MCInst_MC3_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC3_v2_2Inst_1_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC3_v3_0Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_2[2]), .Z(MCInst_MC3_v3_0[1]) );
  XOR2_X1 MCInst_MC3_v3_1Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_1_0_), .Z(MCInst_MC3_v3_1[1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U2 ( .A(MCInst_MC3_v3_3Inst_1_n3), .B(
        MCInst_MC3_v3_2[2]), .ZN(MCInst_MC3_v3_3[1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_1_0_), .ZN(MCInst_MC3_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_3[0]), .Z(MCInst_MC3_v0_0[2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_2_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v0_3[0]), .Z(MCInst_MC3_v0_1[2]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_2_U1 ( .A(MCInst_MC3_v0_0[3]), .B(
        MCInst_MC3_v0_3[0]), .Z(MCInst_MC3_v0_2[2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U2 ( .A(MCInst_MC3_v1_1Inst_2_n3), .B(
        MCInst_MC3_v1_0[3]), .ZN(MCInst_MC3_v1_1[2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U2 ( .A(MCInst_MC3_v1_2Inst_2_n3), .B(
        Red_MCInst_MC3_v1_1_0_), .ZN(MCInst_MC3_v1_2[2]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U2 ( .A(MCInst_MC3_v2_1Inst_2_n3), .B(
        MCInst_MC3_v2_0[0]), .ZN(MCInst_MC3_v2_1[2]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U2 ( .A(MCInst_MC3_v2_2Inst_2_n3), .B(
        MCInst_MC3_v2_0[0]), .ZN(MCInst_MC3_v2_2[2]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC3_v2_3Inst_2_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_3[2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U2 ( .A(MCInst_MC3_v3_1Inst_2_n3), .B(
        MCInst_MC3_v3_2[2]), .ZN(MCInst_MC3_v3_1[2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[2]), .ZN(MCInst_MC3_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC3_v3_3Inst_2_U1 ( .A(MCInst_MC3_v3_0[2]), .B(
        MCInst_MC3_v3_2[2]), .Z(MCInst_MC3_v3_3[2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_3_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_3[0]), .Z(MCInst_MC3_v0_1[3]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_3_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_3[3]), .Z(MCInst_MC3_v0_2[3]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_3_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        Red_MCInst_MC3_v1_1_0_), .Z(MCInst_MC3_v1_1[3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U3 ( .A(MCInst_MC3_v1_2Inst_3_n6), .B(
        MCInst_MC3_v1_2Inst_3_n5), .ZN(MCInst_MC3_v1_2[3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U2 ( .A(Red_MCInst_MC3_v1_1_0_), .B(
        MCInst_MC3_v1_0[3]), .ZN(MCInst_MC3_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC3_v1_2Inst_3_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .Z(MCInst_MC3_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC3_v2_1Inst_3_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[0]), .Z(MCInst_MC3_v2_1[3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U2 ( .A(MCInst_MC3_v2_2Inst_3_n3), .B(
        MCInst_MC3_v2_0[0]), .ZN(MCInst_MC3_v2_2[3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U2 ( .A(MCInst_MC3_v2_3Inst_3_n3), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_3[3]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .ZN(MCInst_MC3_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC3_v3_1Inst_3_U1 ( .A(MCInst_MC3_v3_0[2]), .B(
        Red_MCInst_MC3_v3_1_0_), .Z(MCInst_MC3_v3_1[3]) );
  XOR2_X1 MCInst_MC3_v3_3Inst_3_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_1_0_), .Z(MCInst_MC3_v3_3[3]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_0_n8), .B(MCInst_MC3_r0Inst_XORInst_0_0_n7), .ZN(MC_output[48]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_0[0]), .B(
        MCInst_MC3_v1_0[0]), .ZN(MCInst_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v3_2[2]), .Z(MCInst_MC3_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_1_n8), .B(MCInst_MC3_r0Inst_XORInst_0_1_n7), .ZN(MC_output[49]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_0[1]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_0[1]), .B(
        MCInst_MC3_v3_0[1]), .Z(MCInst_MC3_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_2_n8), .B(MCInst_MC3_r0Inst_XORInst_0_2_n7), .ZN(MC_output[50]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_0[2]), .B(
        Red_MCInst_MC3_v1_1_0_), .ZN(MCInst_MC3_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_0[2]), .B(
        MCInst_MC3_v3_0[2]), .Z(MCInst_MC3_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_3_n8), .B(MCInst_MC3_r0Inst_XORInst_0_3_n7), .ZN(MC_output[51]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        MCInst_MC3_v1_0[3]), .ZN(MCInst_MC3_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_0[3]), .B(
        Red_MCInst_MC3_v3_1_0_), .Z(MCInst_MC3_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_0_n8), .B(MCInst_MC3_r1Inst_XORInst_0_0_n7), .ZN(MC_output[32]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_1[0]), .B(
        MCInst_MC3_v1_1[0]), .ZN(MCInst_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_0[3]), .B(
        MCInst_MC3_v3_1[0]), .Z(MCInst_MC3_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_1_n8), .B(MCInst_MC3_r1Inst_XORInst_0_1_n7), .ZN(MC_output[33]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v1_1[1]), .ZN(MCInst_MC3_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_1[1]), .B(
        MCInst_MC3_v3_1[1]), .Z(MCInst_MC3_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_2_n8), .B(MCInst_MC3_r1Inst_XORInst_0_2_n7), .ZN(MC_output[34]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_1[2]), .B(
        MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_1[2]), .B(
        MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_3_n8), .B(MCInst_MC3_r1Inst_XORInst_0_3_n7), .ZN(MC_output[35]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_1[3]), .B(
        MCInst_MC3_v1_1[3]), .ZN(MCInst_MC3_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_1[3]), .B(
        MCInst_MC3_v3_1[3]), .Z(MCInst_MC3_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_0_n8), .B(MCInst_MC3_r2Inst_XORInst_0_0_n7), .ZN(MC_output[16]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_2[0]), .B(
        MCInst_MC3_v1_2[0]), .ZN(MCInst_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_2[0]), .B(
        MCInst_MC3_v3_2[0]), .Z(MCInst_MC3_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_1_n8), .B(MCInst_MC3_r2Inst_XORInst_0_1_n7), .ZN(MC_output[17]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_2[1]), .B(
        MCInst_MC3_v1_2[1]), .ZN(MCInst_MC3_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_2[1]), .B(
        Red_MCInst_MC3_v3_1_0_), .Z(MCInst_MC3_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_2_n8), .B(MCInst_MC3_r2Inst_XORInst_0_2_n7), .ZN(MC_output[18]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_2[2]), .B(
        MCInst_MC3_v1_2[2]), .ZN(MCInst_MC3_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_2[2]), .Z(MCInst_MC3_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_3_n8), .B(MCInst_MC3_r2Inst_XORInst_0_3_n7), .ZN(MC_output[19]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_2[3]), .B(
        MCInst_MC3_v1_2[3]), .ZN(MCInst_MC3_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_2[3]), .B(
        MCInst_MC3_v3_2[3]), .Z(MCInst_MC3_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_0_n8), .B(MCInst_MC3_r3Inst_XORInst_0_0_n7), .ZN(MC_output[0]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_3[0]), .B(
        MCInst_MC3_v1_0[3]), .ZN(MCInst_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_3[0]), .B(
        MCInst_MC3_v3_3[0]), .Z(MCInst_MC3_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_1_n8), .B(MCInst_MC3_r3Inst_XORInst_0_1_n7), .ZN(MC_output[1]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v1_3[1]), .ZN(MCInst_MC3_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_3[1]), .B(
        MCInst_MC3_v3_3[1]), .Z(MCInst_MC3_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_2_n8), .B(MCInst_MC3_r3Inst_XORInst_0_2_n7), .ZN(MC_output[2]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_3[2]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_0[3]), .B(
        MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_3_n8), .B(MCInst_MC3_r3Inst_XORInst_0_3_n7), .ZN(MC_output[3]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_3[3]), .B(
        Red_MCInst_MC3_v1_1_0_), .ZN(MCInst_MC3_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v3_3[3]), .Z(MCInst_MC3_r3Inst_XORInst_0_3_n8) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(MC_output[0]), .CK(clk), .Q(
        SubCellInput2[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(MC_output[1]), .CK(clk), .Q(
        SubCellInput2[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(MC_output[2]), .CK(clk), .Q(
        SubCellInput2[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(MC_output[3]), .CK(clk), .Q(
        SubCellInput2[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(MC_output[4]), .CK(clk), .Q(
        SubCellInput2[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(MC_output[5]), .CK(clk), .Q(
        SubCellInput2[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(MC_output[6]), .CK(clk), .Q(
        SubCellInput2[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(MC_output[7]), .CK(clk), .Q(
        SubCellInput2[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(MC_output[8]), .CK(clk), .Q(
        SubCellInput2[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(MC_output[9]), .CK(clk), .Q(
        SubCellInput2[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(MC_output[10]), .CK(clk), .Q(
        SubCellInput2[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(MC_output[11]), .CK(clk), .Q(
        SubCellInput2[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(MC_output[12]), .CK(clk), .Q(
        SubCellInput2[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(MC_output[13]), .CK(clk), .Q(
        SubCellInput2[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(MC_output[14]), .CK(clk), .Q(
        SubCellInput2[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(MC_output[15]), .CK(clk), .Q(
        SubCellInput2[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(MC_output[16]), .CK(clk), .Q(
        SubCellInput2[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(MC_output[17]), .CK(clk), .Q(
        SubCellInput2[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(MC_output[18]), .CK(clk), .Q(
        SubCellInput2[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(MC_output[19]), .CK(clk), .Q(
        SubCellInput2[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(MC_output[20]), .CK(clk), .Q(
        SubCellInput2[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(MC_output[21]), .CK(clk), .Q(
        SubCellInput2[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(MC_output[22]), .CK(clk), .Q(
        SubCellInput2[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(MC_output[23]), .CK(clk), .Q(
        SubCellInput2[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(MC_output[24]), .CK(clk), .Q(
        SubCellInput2[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(MC_output[25]), .CK(clk), .Q(
        SubCellInput2[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(MC_output[26]), .CK(clk), .Q(
        SubCellInput2[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(MC_output[27]), .CK(clk), .Q(
        SubCellInput2[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(MC_output[28]), .CK(clk), .Q(
        SubCellInput2[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(MC_output[29]), .CK(clk), .Q(
        SubCellInput2[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(MC_output[30]), .CK(clk), .Q(
        SubCellInput2[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(MC_output[31]), .CK(clk), .Q(
        SubCellInput2[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(MC_output[32]), .CK(clk), .Q(
        SubCellInput2[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(MC_output[33]), .CK(clk), .Q(
        SubCellInput2[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(MC_output[34]), .CK(clk), .Q(
        SubCellInput2[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(MC_output[35]), .CK(clk), .Q(
        SubCellInput2[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(MC_output[36]), .CK(clk), .Q(
        SubCellInput2[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(MC_output[37]), .CK(clk), .Q(
        SubCellInput2[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(MC_output[38]), .CK(clk), .Q(
        SubCellInput2[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(MC_output[39]), .CK(clk), .Q(
        SubCellInput2[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(MC_output[40]), .CK(clk), .Q(
        SubCellInput2[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(MC_output[41]), .CK(clk), .Q(
        SubCellInput2[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(MC_output[42]), .CK(clk), .Q(
        SubCellInput2[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(MC_output[43]), .CK(clk), .Q(
        SubCellInput2[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(MC_output[44]), .CK(clk), .Q(
        SubCellInput2[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(MC_output[45]), .CK(clk), .Q(
        SubCellInput2[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(MC_output[46]), .CK(clk), .Q(
        SubCellInput2[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(MC_output[47]), .CK(clk), .Q(
        SubCellInput2[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(MC_output[48]), .CK(clk), .Q(
        SubCellInput2[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(MC_output[49]), .CK(clk), .Q(
        SubCellInput2[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(MC_output[50]), .CK(clk), .Q(
        SubCellInput2[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(MC_output[51]), .CK(clk), .Q(
        SubCellInput2[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(MC_output[52]), .CK(clk), .Q(
        SubCellInput2[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(MC_output[53]), .CK(clk), .Q(
        SubCellInput2[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(MC_output[54]), .CK(clk), .Q(
        SubCellInput2[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(MC_output[55]), .CK(clk), .Q(
        SubCellInput2[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(MC_output[56]), .CK(clk), .Q(
        SubCellInput2[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(MC_output[57]), .CK(clk), .Q(
        SubCellInput2[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(MC_output[58]), .CK(clk), .Q(
        SubCellInput2[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(MC_output[59]), .CK(clk), .Q(
        SubCellInput2[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(MC_output[60]), .CK(clk), .Q(
        SubCellInput2[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(MC_output[61]), .CK(clk), .Q(
        SubCellInput2[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(MC_output[62]), .CK(clk), .Q(
        SubCellInput2[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(MC_output[63]), .CK(clk), .Q(
        SubCellInput2[63]), .QN() );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_0_U4 ( .A1(SubCellInput2[2]), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_0_U3 ( .A(SubCellInput2[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U2 ( .A(SubCellInput2[0]), .B(
        SubCellInput2[3]), .ZN(SubCellInst2_LFInst_0_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_0_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_0_LFInst_0_n5), .B(
        SubCellInst2_LFInst_0_LFInst_0_n7), .Z(MCInst2_MC0_v3_2[3]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n25), .ZN(MCInst2_MC0_v3_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_1_U8 ( .A1(SubCellInput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_1_U7 ( .A(SubCellInput2[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n21), .A2(SubCellInput2[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U4 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U2 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_1_U1 ( .A(SubCellInput2[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n28), .ZN(Red_MCInst2_MC0_v3_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_2_U6 ( .A(SubCellInput2[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_0_LFInst_2_n25), .B(SubCellInput2[2]), .Z(
        SubCellInst2_LFInst_0_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U4 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n23), .A2(SubCellInput2[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_0_LFInst_2_n22), .B(SubCellInput2[1]), .Z(
        SubCellInst2_LFInst_0_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_2_U1 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U9 ( .A1(SubCellInput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n23), .A2(SubCellInput2[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_3_U7 ( .A1(SubCellInput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U4 ( .A1(SubCellInput2[2]), .A2(
        SubCellInput2[0]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_3_U3 ( .A(SubCellInput2[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U2 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n25), .ZN(MCInst2_MC0_v3_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_0_U4 ( .A1(SubCellInput2[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_0_U3 ( .A(SubCellInput2[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U2 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[7]), .ZN(SubCellInst2_LFInst_1_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_1_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_1_LFInst_0_n5), .B(
        SubCellInst2_LFInst_1_LFInst_0_n7), .Z(MCInst2_MC3_v3_2[3]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n25), .ZN(MCInst2_MC3_v3_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_1_U8 ( .A1(SubCellInput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_1_U7 ( .A(SubCellInput2[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n21), .A2(SubCellInput2[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U4 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U2 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_1_U1 ( .A(SubCellInput2[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n28), .ZN(Red_MCInst2_MC3_v3_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_2_U6 ( .A(SubCellInput2[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_1_LFInst_2_n25), .B(SubCellInput2[6]), .Z(
        SubCellInst2_LFInst_1_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U4 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n23), .A2(SubCellInput2[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_1_LFInst_2_n22), .B(SubCellInput2[5]), .Z(
        SubCellInst2_LFInst_1_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_2_U1 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U9 ( .A1(SubCellInput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n23), .A2(SubCellInput2[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_3_U7 ( .A1(SubCellInput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U4 ( .A1(SubCellInput2[6]), .A2(
        SubCellInput2[4]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_3_U3 ( .A(SubCellInput2[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U2 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n25), .ZN(MCInst2_MC3_v3_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_0_U4 ( .A1(SubCellInput2[10]), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_0_U3 ( .A(SubCellInput2[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U2 ( .A(SubCellInput2[8]), .B(
        SubCellInput2[11]), .ZN(SubCellInst2_LFInst_2_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_2_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_2_LFInst_0_n5), .B(
        SubCellInst2_LFInst_2_LFInst_0_n7), .Z(MCInst2_MC2_v3_2[3]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n25), .ZN(MCInst2_MC2_v3_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_1_U8 ( .A1(SubCellInput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_1_U7 ( .A(SubCellInput2[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n21), .A2(SubCellInput2[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U4 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U2 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_1_U1 ( .A(SubCellInput2[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n28), .ZN(Red_MCInst2_MC2_v3_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_2_U6 ( .A(SubCellInput2[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_2_LFInst_2_n25), .B(SubCellInput2[10]), .Z(
        SubCellInst2_LFInst_2_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U4 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n23), .A2(SubCellInput2[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_2_LFInst_2_n22), .B(SubCellInput2[9]), .Z(
        SubCellInst2_LFInst_2_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_2_U1 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U9 ( .A1(SubCellInput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n23), .A2(SubCellInput2[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_3_U7 ( .A1(SubCellInput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U4 ( .A1(SubCellInput2[10]), .A2(
        SubCellInput2[8]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_3_U3 ( .A(SubCellInput2[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U2 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n25), .ZN(MCInst2_MC2_v3_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_0_U4 ( .A1(SubCellInput2[14]), .A2(
        SubCellInst2_LFInst_3_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_0_U3 ( .A(SubCellInput2[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U2 ( .A(SubCellInput2[12]), .B(
        SubCellInput2[15]), .ZN(SubCellInst2_LFInst_3_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_3_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_3_LFInst_0_n5), .B(
        SubCellInst2_LFInst_3_LFInst_0_n7), .Z(MCInst2_MC1_v3_2[3]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n25), .ZN(MCInst2_MC1_v3_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_1_U8 ( .A1(SubCellInput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_1_U7 ( .A(SubCellInput2[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n21), .A2(SubCellInput2[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U4 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U2 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_1_U1 ( .A(SubCellInput2[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n28), .ZN(Red_MCInst2_MC1_v3_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_2_U6 ( .A(SubCellInput2[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_3_LFInst_2_n25), .B(SubCellInput2[14]), .Z(
        SubCellInst2_LFInst_3_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U4 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n23), .A2(SubCellInput2[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_3_LFInst_2_n22), .B(SubCellInput2[13]), .Z(
        SubCellInst2_LFInst_3_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_2_U1 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U9 ( .A1(SubCellInput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n23), .A2(SubCellInput2[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_3_U7 ( .A1(SubCellInput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U4 ( .A1(SubCellInput2[14]), .A2(
        SubCellInput2[12]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_3_U3 ( .A(SubCellInput2[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U2 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n25), .ZN(MCInst2_MC1_v3_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_0_U4 ( .A1(SubCellInput2[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_0_U3 ( .A(SubCellInput2[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U2 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[19]), .ZN(SubCellInst2_LFInst_4_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_4_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_4_LFInst_0_n5), .B(
        SubCellInst2_LFInst_4_LFInst_0_n7), .Z(MCInst2_MC1_v2_3[1]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n25), .ZN(MCInst2_MC1_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_1_U8 ( .A1(SubCellInput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_1_U7 ( .A(SubCellInput2[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n21), .A2(SubCellInput2[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U4 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U2 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_1_U1 ( .A(SubCellInput2[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n28), .ZN(MCInst2_MC1_v2_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U8 ( .A1(SubCellInput2[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U7 ( .A1(SubCellInput2[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_2_U6 ( .A(SubCellInput2[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_4_LFInst_2_n23), .B(SubCellInput2[18]), .Z(
        SubCellInst2_LFInst_4_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U3 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n22), .A2(SubCellInput2[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U1 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U9 ( .A1(SubCellInput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n23), .A2(SubCellInput2[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_4_LFInst_3_U7 ( .A1(SubCellInput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U4 ( .A1(SubCellInput2[18]), .A2(
        SubCellInput2[16]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_3_U3 ( .A(SubCellInput2[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U2 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n25), .ZN(MCInst2_MC1_v2_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_0_U4 ( .A1(SubCellInput2[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_0_U3 ( .A(SubCellInput2[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U2 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[23]), .ZN(SubCellInst2_LFInst_5_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_5_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_5_LFInst_0_n5), .B(
        SubCellInst2_LFInst_5_LFInst_0_n7), .Z(MCInst2_MC0_v2_3[1]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n25), .ZN(MCInst2_MC0_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_1_U8 ( .A1(SubCellInput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_1_U7 ( .A(SubCellInput2[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n21), .A2(SubCellInput2[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U4 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U2 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_1_U1 ( .A(SubCellInput2[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n28), .ZN(MCInst2_MC0_v2_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U8 ( .A1(SubCellInput2[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U7 ( .A1(SubCellInput2[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_2_U6 ( .A(SubCellInput2[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_5_LFInst_2_n23), .B(SubCellInput2[22]), .Z(
        SubCellInst2_LFInst_5_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U3 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n22), .A2(SubCellInput2[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U1 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U9 ( .A1(SubCellInput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n23), .A2(SubCellInput2[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_5_LFInst_3_U7 ( .A1(SubCellInput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U4 ( .A1(SubCellInput2[22]), .A2(
        SubCellInput2[20]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_3_U3 ( .A(SubCellInput2[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U2 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n25), .ZN(MCInst2_MC0_v2_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_0_U4 ( .A1(SubCellInput2[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_0_U3 ( .A(SubCellInput2[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U2 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[27]), .ZN(SubCellInst2_LFInst_6_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_6_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_6_LFInst_0_n5), .B(
        SubCellInst2_LFInst_6_LFInst_0_n7), .Z(MCInst2_MC3_v2_3[1]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n25), .ZN(MCInst2_MC3_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_1_U8 ( .A1(SubCellInput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_1_U7 ( .A(SubCellInput2[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n21), .A2(SubCellInput2[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U4 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U2 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_1_U1 ( .A(SubCellInput2[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n28), .ZN(MCInst2_MC3_v2_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U8 ( .A1(SubCellInput2[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U7 ( .A1(SubCellInput2[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_2_U6 ( .A(SubCellInput2[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_6_LFInst_2_n23), .B(SubCellInput2[26]), .Z(
        SubCellInst2_LFInst_6_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U3 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n22), .A2(SubCellInput2[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U1 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U9 ( .A1(SubCellInput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n23), .A2(SubCellInput2[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_6_LFInst_3_U7 ( .A1(SubCellInput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U4 ( .A1(SubCellInput2[26]), .A2(
        SubCellInput2[24]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_3_U3 ( .A(SubCellInput2[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U2 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n25), .ZN(MCInst2_MC3_v2_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_0_U4 ( .A1(SubCellInput2[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_0_U3 ( .A(SubCellInput2[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U2 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[31]), .ZN(SubCellInst2_LFInst_7_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_7_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_7_LFInst_0_n5), .B(
        SubCellInst2_LFInst_7_LFInst_0_n7), .Z(MCInst2_MC2_v2_3[1]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n25), .ZN(MCInst2_MC2_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_1_U8 ( .A1(SubCellInput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_1_U7 ( .A(SubCellInput2[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n21), .A2(SubCellInput2[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U4 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U2 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_1_U1 ( .A(SubCellInput2[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n28), .ZN(MCInst2_MC2_v2_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U8 ( .A1(SubCellInput2[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U7 ( .A1(SubCellInput2[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_2_U6 ( .A(SubCellInput2[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_7_LFInst_2_n23), .B(SubCellInput2[30]), .Z(
        SubCellInst2_LFInst_7_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U3 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n22), .A2(SubCellInput2[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U1 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U9 ( .A1(SubCellInput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n23), .A2(SubCellInput2[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_7_LFInst_3_U7 ( .A1(SubCellInput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U4 ( .A1(SubCellInput2[30]), .A2(
        SubCellInput2[28]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_3_U3 ( .A(SubCellInput2[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U2 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n25), .ZN(MCInst2_MC2_v2_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_0_U4 ( .A1(SubCellInput2[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_0_U3 ( .A(SubCellInput2[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U2 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[35]), .ZN(SubCellInst2_LFInst_8_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_8_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_8_LFInst_0_n5), .B(
        SubCellInst2_LFInst_8_LFInst_0_n7), .Z(MCInst2_MC2_v1_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n25), .ZN(MCInst2_MC2_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_1_U8 ( .A1(SubCellInput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_1_U7 ( .A(SubCellInput2[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n21), .A2(SubCellInput2[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U4 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U2 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_1_U1 ( .A(SubCellInput2[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U9 ( .A1(SubCellInput2[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U8 ( .A1(SubCellInput2[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_2_U7 ( .A(SubCellInput2[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_8_LFInst_2_n23), .B(SubCellInput2[34]), .Z(
        SubCellInst2_LFInst_8_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U4 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n22), .A2(SubCellInput2[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U2 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n28), .ZN(Red_MCInst2_MC2_v1_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n25), .ZN(MCInst2_MC2_v1_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U8 ( .A1(SubCellInput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n23), .A2(SubCellInput2[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_3_U6 ( .A1(SubCellInput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U3 ( .A1(SubCellInput2[34]), .A2(
        SubCellInput2[32]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_3_U2 ( .A(SubCellInput2[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U1 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_0_U4 ( .A1(SubCellInput2[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_0_U3 ( .A(SubCellInput2[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U2 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[39]), .ZN(SubCellInst2_LFInst_9_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_9_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_9_LFInst_0_n5), .B(
        SubCellInst2_LFInst_9_LFInst_0_n7), .Z(MCInst2_MC1_v1_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n25), .ZN(MCInst2_MC1_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_1_U8 ( .A1(SubCellInput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_1_U7 ( .A(SubCellInput2[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n21), .A2(SubCellInput2[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U4 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U2 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_1_U1 ( .A(SubCellInput2[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U9 ( .A1(SubCellInput2[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U8 ( .A1(SubCellInput2[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_2_U7 ( .A(SubCellInput2[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_9_LFInst_2_n23), .B(SubCellInput2[38]), .Z(
        SubCellInst2_LFInst_9_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U4 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n22), .A2(SubCellInput2[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U2 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n28), .ZN(Red_MCInst2_MC1_v1_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n25), .ZN(MCInst2_MC1_v1_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U8 ( .A1(SubCellInput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n23), .A2(SubCellInput2[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_3_U6 ( .A1(SubCellInput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U3 ( .A1(SubCellInput2[38]), .A2(
        SubCellInput2[36]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_3_U2 ( .A(SubCellInput2[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U1 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_0_U4 ( .A1(SubCellInput2[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_0_U3 ( .A(SubCellInput2[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U2 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[43]), .ZN(SubCellInst2_LFInst_10_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_10_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_10_LFInst_0_n5), .B(
        SubCellInst2_LFInst_10_LFInst_0_n7), .Z(MCInst2_MC0_v1_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n25), .ZN(MCInst2_MC0_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_1_U8 ( .A1(SubCellInput2[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_1_U7 ( .A(SubCellInput2[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n21), .A2(SubCellInput2[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U4 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U2 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_1_U1 ( .A(SubCellInput2[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U9 ( .A1(SubCellInput2[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U8 ( .A1(SubCellInput2[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_2_U7 ( .A(SubCellInput2[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_10_LFInst_2_n23), .B(SubCellInput2[42]), .Z(
        SubCellInst2_LFInst_10_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U4 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n22), .A2(SubCellInput2[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U2 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n28), .ZN(Red_MCInst2_MC0_v1_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n25), .ZN(MCInst2_MC0_v1_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U8 ( .A1(SubCellInput2[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n23), .A2(SubCellInput2[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_3_U6 ( .A1(SubCellInput2[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U3 ( .A1(SubCellInput2[42]), .A2(
        SubCellInput2[40]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_3_U2 ( .A(SubCellInput2[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U1 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_0_U4 ( .A1(SubCellInput2[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_0_U3 ( .A(SubCellInput2[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U2 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[47]), .ZN(SubCellInst2_LFInst_11_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_11_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_11_LFInst_0_n5), .B(
        SubCellInst2_LFInst_11_LFInst_0_n7), .Z(MCInst2_MC3_v1_0[0]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n25), .ZN(MCInst2_MC3_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_1_U8 ( .A1(SubCellInput2[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_1_U7 ( .A(SubCellInput2[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n21), .A2(SubCellInput2[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U4 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U2 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_1_U1 ( .A(SubCellInput2[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U9 ( .A1(SubCellInput2[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U8 ( .A1(SubCellInput2[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_2_U7 ( .A(SubCellInput2[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_11_LFInst_2_n23), .B(SubCellInput2[46]), .Z(
        SubCellInst2_LFInst_11_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U4 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n22), .A2(SubCellInput2[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U2 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n28), .ZN(Red_MCInst2_MC3_v1_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n25), .ZN(MCInst2_MC3_v1_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U8 ( .A1(SubCellInput2[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n23), .A2(SubCellInput2[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_3_U6 ( .A1(SubCellInput2[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U3 ( .A1(SubCellInput2[46]), .A2(
        SubCellInput2[44]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_3_U2 ( .A(SubCellInput2[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U1 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_0_U4 ( .A1(SubCellInput2[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_0_U3 ( .A(SubCellInput2[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U2 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[51]), .ZN(SubCellInst2_LFInst_12_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_12_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_12_LFInst_0_n5), .B(
        SubCellInst2_LFInst_12_LFInst_0_n7), .Z(Red_MCInst2_MC3_v0_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n25), .ZN(MCInst2_MC3_v0_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_1_U8 ( .A1(SubCellInput2[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_1_U7 ( .A(SubCellInput2[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n21), .A2(SubCellInput2[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U4 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U2 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_1_U1 ( .A(SubCellInput2[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n28), .ZN(MCInst2_MC3_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U8 ( .A1(SubCellInput2[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U7 ( .A1(SubCellInput2[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_2_U6 ( .A(SubCellInput2[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_12_LFInst_2_n23), .B(SubCellInput2[50]), .Z(
        SubCellInst2_LFInst_12_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U3 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n22), .A2(SubCellInput2[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U1 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U9 ( .A1(SubCellInput2[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n23), .A2(SubCellInput2[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_3_U7 ( .A1(SubCellInput2[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U4 ( .A1(SubCellInput2[50]), .A2(
        SubCellInput2[48]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_3_U3 ( .A(SubCellInput2[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U2 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n25), .ZN(MCInst2_MC3_v0_3[0]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_0_U4 ( .A1(SubCellInput2[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_0_U3 ( .A(SubCellInput2[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U2 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[55]), .ZN(SubCellInst2_LFInst_13_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_13_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_13_LFInst_0_n5), .B(
        SubCellInst2_LFInst_13_LFInst_0_n7), .Z(Red_MCInst2_MC2_v0_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n25), .ZN(MCInst2_MC2_v0_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_1_U8 ( .A1(SubCellInput2[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_1_U7 ( .A(SubCellInput2[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n21), .A2(SubCellInput2[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U4 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U2 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_1_U1 ( .A(SubCellInput2[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n28), .ZN(MCInst2_MC2_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U8 ( .A1(SubCellInput2[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U7 ( .A1(SubCellInput2[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_2_U6 ( .A(SubCellInput2[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_13_LFInst_2_n23), .B(SubCellInput2[54]), .Z(
        SubCellInst2_LFInst_13_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U3 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n22), .A2(SubCellInput2[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U1 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U9 ( .A1(SubCellInput2[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n23), .A2(SubCellInput2[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_3_U7 ( .A1(SubCellInput2[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U4 ( .A1(SubCellInput2[54]), .A2(
        SubCellInput2[52]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_3_U3 ( .A(SubCellInput2[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U2 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n25), .ZN(MCInst2_MC2_v0_3[0]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_0_U4 ( .A1(SubCellInput2[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_0_U3 ( .A(SubCellInput2[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U2 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[59]), .ZN(SubCellInst2_LFInst_14_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_14_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_14_LFInst_0_n5), .B(
        SubCellInst2_LFInst_14_LFInst_0_n7), .Z(Red_MCInst2_MC1_v0_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n25), .ZN(MCInst2_MC1_v0_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_1_U8 ( .A1(SubCellInput2[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_1_U7 ( .A(SubCellInput2[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n21), .A2(SubCellInput2[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U4 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U2 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_1_U1 ( .A(SubCellInput2[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n28), .ZN(MCInst2_MC1_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U8 ( .A1(SubCellInput2[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U7 ( .A1(SubCellInput2[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_2_U6 ( .A(SubCellInput2[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_14_LFInst_2_n23), .B(SubCellInput2[58]), .Z(
        SubCellInst2_LFInst_14_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U3 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n22), .A2(SubCellInput2[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U1 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U9 ( .A1(SubCellInput2[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n23), .A2(SubCellInput2[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_3_U7 ( .A1(SubCellInput2[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U4 ( .A1(SubCellInput2[58]), .A2(
        SubCellInput2[56]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_3_U3 ( .A(SubCellInput2[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U2 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n25), .ZN(MCInst2_MC1_v0_3[0]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_0_U4 ( .A1(SubCellInput2[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_0_n6), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_0_U3 ( .A(SubCellInput2[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n6) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U2 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[63]), .ZN(SubCellInst2_LFInst_15_LFInst_0_n5) );
  XOR2_X2 SubCellInst2_LFInst_15_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_15_LFInst_0_n5), .B(
        SubCellInst2_LFInst_15_LFInst_0_n7), .Z(Red_MCInst2_MC0_v0_1_0_) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n25), .ZN(MCInst2_MC0_v0_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_1_U8 ( .A1(SubCellInput2[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_1_U7 ( .A(SubCellInput2[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n21), .A2(SubCellInput2[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U4 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U2 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_1_U1 ( .A(SubCellInput2[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U9 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n28), .ZN(MCInst2_MC0_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U8 ( .A1(SubCellInput2[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U7 ( .A1(SubCellInput2[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_2_U6 ( .A(SubCellInput2[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U5 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U4 ( .A(
        SubCellInst2_LFInst_15_LFInst_2_n23), .B(SubCellInput2[62]), .Z(
        SubCellInst2_LFInst_15_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U3 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U2 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n22), .A2(SubCellInput2[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U1 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U9 ( .A1(SubCellInput2[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n23), .A2(SubCellInput2[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_3_U7 ( .A1(SubCellInput2[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U4 ( .A1(SubCellInput2[62]), .A2(
        SubCellInput2[60]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_3_U3 ( .A(SubCellInput2[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U2 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n25), .ZN(MCInst2_MC0_v0_3[0]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U2 ( .A(MCInst2_MC0_v0_2Inst_0_n3), .B(
        MCInst2_MC0_v0_3[0]), .ZN(MCInst2_MC0_v0_2[0]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_0[3]), .ZN(MCInst2_MC0_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_0_U1 ( .A(Red_MCInst2_MC0_v1_1_0_), .B(
        MCInst2_MC0_v1_0[3]), .Z(MCInst2_MC0_v1_1[0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U2 ( .A(MCInst2_MC0_v1_2Inst_0_n3), .B(
        MCInst2_MC0_v1_0[3]), .ZN(MCInst2_MC0_v1_2[0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U1 ( .A(MCInst2_MC0_v1_3[2]), .B(
        Red_MCInst2_MC0_v1_1_0_), .ZN(MCInst2_MC0_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_0_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[3]), .Z(MCInst2_MC0_v2_1[0]) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_0_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[0]), .Z(MCInst2_MC0_v2_2[0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U3 ( .A(MCInst2_MC0_v2_3Inst_0_n6), .B(
        MCInst2_MC0_v2_3Inst_0_n5), .ZN(MCInst2_MC0_v2_3[0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        MCInst2_MC0_v2_0[0]), .ZN(MCInst2_MC0_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_0_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(MCInst2_MC0_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_0_U1 ( .A(Red_MCInst2_MC0_v3_1_0_), .B(
        MCInst2_MC0_v3_2[2]), .Z(MCInst2_MC0_v3_1[0]) );
  XOR2_X1 MCInst2_MC0_v3_2Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[2]), .Z(MCInst2_MC0_v3_2[0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U2 ( .A(MCInst2_MC0_v3_3Inst_0_n3), .B(
        MCInst2_MC0_v3_2[2]), .ZN(MCInst2_MC0_v3_3[0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[2]), .ZN(MCInst2_MC0_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_1_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        MCInst2_MC0_v0_3[0]), .Z(MCInst2_MC0_v0_0[1]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_1_U1 ( .A(MCInst2_MC0_v0_0[3]), .B(
        MCInst2_MC0_v0_3[3]), .Z(MCInst2_MC0_v0_1[1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U2 ( .A(MCInst2_MC0_v0_2Inst_1_n3), .B(
        MCInst2_MC0_v0_3[0]), .ZN(MCInst2_MC0_v0_2[1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_3[3]), .ZN(MCInst2_MC0_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_3[0]), .Z(MCInst2_MC0_v0_3[1]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_1_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        Red_MCInst2_MC0_v1_1_0_), .Z(MCInst2_MC0_v1_1[1]) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_1_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .Z(MCInst2_MC0_v1_2[1]) );
  XOR2_X1 MCInst2_MC0_v1_3Inst_1_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_0[3]), .Z(MCInst2_MC0_v1_3[1]) );
  XOR2_X1 MCInst2_MC0_v2_0Inst_1_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[0]), .Z(MCInst2_MC0_v2_0[1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U2 ( .A(MCInst2_MC0_v2_1Inst_1_n3), .B(
        MCInst2_MC0_v2_0[0]), .ZN(MCInst2_MC0_v2_1[1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U3 ( .A(MCInst2_MC0_v2_2Inst_1_n6), .B(
        MCInst2_MC0_v2_2Inst_1_n5), .ZN(MCInst2_MC0_v2_2[1]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        MCInst2_MC0_v2_0[0]), .ZN(MCInst2_MC0_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_1_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(MCInst2_MC0_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC0_v3_0Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_2[2]), .Z(MCInst2_MC0_v3_0[1]) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_1_0_), .Z(MCInst2_MC0_v3_1[1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U2 ( .A(MCInst2_MC0_v3_3Inst_1_n3), .B(
        MCInst2_MC0_v3_2[2]), .ZN(MCInst2_MC0_v3_3[1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_1_0_), .ZN(MCInst2_MC0_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_3[0]), .Z(MCInst2_MC0_v0_0[2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_2_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        MCInst2_MC0_v0_3[0]), .Z(MCInst2_MC0_v0_1[2]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_2_U1 ( .A(MCInst2_MC0_v0_0[3]), .B(
        MCInst2_MC0_v0_3[0]), .Z(MCInst2_MC0_v0_2[2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U2 ( .A(MCInst2_MC0_v1_1Inst_2_n3), .B(
        MCInst2_MC0_v1_0[3]), .ZN(MCInst2_MC0_v1_1[2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U2 ( .A(MCInst2_MC0_v1_2Inst_2_n3), .B(
        Red_MCInst2_MC0_v1_1_0_), .ZN(MCInst2_MC0_v1_2[2]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U2 ( .A(MCInst2_MC0_v2_1Inst_2_n3), .B(
        MCInst2_MC0_v2_0[0]), .ZN(MCInst2_MC0_v2_1[2]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U2 ( .A(MCInst2_MC0_v2_2Inst_2_n3), .B(
        MCInst2_MC0_v2_0[0]), .ZN(MCInst2_MC0_v2_2[2]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_2_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(MCInst2_MC0_v2_3[2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U2 ( .A(MCInst2_MC0_v3_1Inst_2_n3), .B(
        MCInst2_MC0_v3_2[2]), .ZN(MCInst2_MC0_v3_1[2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[2]), .ZN(MCInst2_MC0_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_2_U1 ( .A(MCInst2_MC0_v3_0[2]), .B(
        MCInst2_MC0_v3_2[2]), .Z(MCInst2_MC0_v3_3[2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_3[0]), .Z(MCInst2_MC0_v0_1[3]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_3[3]), .Z(MCInst2_MC0_v0_2[3]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_3_U1 ( .A(MCInst2_MC0_v1_3[2]), .B(
        Red_MCInst2_MC0_v1_1_0_), .Z(MCInst2_MC0_v1_1[3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U3 ( .A(MCInst2_MC0_v1_2Inst_3_n6), .B(
        MCInst2_MC0_v1_2Inst_3_n5), .ZN(MCInst2_MC0_v1_2[3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U2 ( .A(Red_MCInst2_MC0_v1_1_0_), .B(
        MCInst2_MC0_v1_0[3]), .ZN(MCInst2_MC0_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_3_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .Z(MCInst2_MC0_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_3_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[0]), .Z(MCInst2_MC0_v2_1[3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U2 ( .A(MCInst2_MC0_v2_2Inst_3_n3), .B(
        MCInst2_MC0_v2_0[0]), .ZN(MCInst2_MC0_v2_2[3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U2 ( .A(MCInst2_MC0_v2_3Inst_3_n3), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_3[3]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .ZN(MCInst2_MC0_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_3_U1 ( .A(MCInst2_MC0_v3_0[2]), .B(
        Red_MCInst2_MC0_v3_1_0_), .Z(MCInst2_MC0_v3_1[3]) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_3_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_1_0_), .Z(MCInst2_MC0_v3_3[3]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[60]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_0[0]), .B(
        MCInst2_MC0_v1_0[0]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        MCInst2_MC0_v3_2[2]), .Z(MCInst2_MC0_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[61]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_0[1]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_0[1]), .B(
        MCInst2_MC0_v3_0[1]), .Z(MCInst2_MC0_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[62]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_0[2]), .B(
        Red_MCInst2_MC0_v1_1_0_), .ZN(MCInst2_MC0_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_0[2]), .B(
        MCInst2_MC0_v3_0[2]), .Z(MCInst2_MC0_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[63]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        MCInst2_MC0_v1_0[3]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_0[3]), .B(
        Red_MCInst2_MC0_v3_1_0_), .Z(MCInst2_MC0_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[44]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_1[0]), .B(
        MCInst2_MC0_v1_1[0]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U1 ( .A(MCInst2_MC0_v0_0[3]), .B(
        MCInst2_MC0_v3_1[0]), .Z(MCInst2_MC0_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[45]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v1_1[1]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_1[1]), .B(
        MCInst2_MC0_v3_1[1]), .Z(MCInst2_MC0_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[46]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_1[2]), .B(
        MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_1[2]), .B(
        MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[47]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_1[3]), .B(
        MCInst2_MC0_v1_1[3]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_1[3]), .B(
        MCInst2_MC0_v3_1[3]), .Z(MCInst2_MC0_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[28]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_2[0]), .B(
        MCInst2_MC0_v1_2[0]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC0_v0_2[0]), .B(
        MCInst2_MC0_v3_2[0]), .Z(MCInst2_MC0_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[29]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_2[1]), .B(
        MCInst2_MC0_v1_2[1]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_2[1]), .B(
        Red_MCInst2_MC0_v3_1_0_), .Z(MCInst2_MC0_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[30]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_2[2]), .B(
        MCInst2_MC0_v1_2[2]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_2[2]), .B(
        MCInst2_MC0_v3_2[2]), .Z(MCInst2_MC0_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[31]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_2[3]), .B(
        MCInst2_MC0_v1_2[3]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_2[3]), .B(
        MCInst2_MC0_v3_2[3]), .Z(MCInst2_MC0_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[12]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_3[0]), .B(
        MCInst2_MC0_v1_0[3]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U1 ( .A(MCInst2_MC0_v0_3[0]), .B(
        MCInst2_MC0_v3_3[0]), .Z(MCInst2_MC0_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[13]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v1_3[1]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_3[1]), .B(
        MCInst2_MC0_v3_3[1]), .Z(MCInst2_MC0_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[14]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_3[2]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_0[3]), .B(
        MCInst2_MC0_v3_3[2]), .Z(MCInst2_MC0_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[15]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_3[3]), .B(
        Red_MCInst2_MC0_v1_1_0_), .ZN(MCInst2_MC0_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        MCInst2_MC0_v3_3[3]), .Z(MCInst2_MC0_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U2 ( .A(MCInst2_MC1_v0_2Inst_0_n3), .B(
        MCInst2_MC1_v0_3[0]), .ZN(MCInst2_MC1_v0_2[0]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_0[3]), .ZN(MCInst2_MC1_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_0_U1 ( .A(Red_MCInst2_MC1_v1_1_0_), .B(
        MCInst2_MC1_v1_0[3]), .Z(MCInst2_MC1_v1_1[0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U2 ( .A(MCInst2_MC1_v1_2Inst_0_n3), .B(
        MCInst2_MC1_v1_0[3]), .ZN(MCInst2_MC1_v1_2[0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U1 ( .A(MCInst2_MC1_v1_3[2]), .B(
        Red_MCInst2_MC1_v1_1_0_), .ZN(MCInst2_MC1_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_0_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[3]), .Z(MCInst2_MC1_v2_1[0]) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_0_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[0]), .Z(MCInst2_MC1_v2_2[0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U3 ( .A(MCInst2_MC1_v2_3Inst_0_n6), .B(
        MCInst2_MC1_v2_3Inst_0_n5), .ZN(MCInst2_MC1_v2_3[0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        MCInst2_MC1_v2_0[0]), .ZN(MCInst2_MC1_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_0_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(MCInst2_MC1_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_0_U1 ( .A(Red_MCInst2_MC1_v3_1_0_), .B(
        MCInst2_MC1_v3_2[2]), .Z(MCInst2_MC1_v3_1[0]) );
  XOR2_X1 MCInst2_MC1_v3_2Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[2]), .Z(MCInst2_MC1_v3_2[0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U2 ( .A(MCInst2_MC1_v3_3Inst_0_n3), .B(
        MCInst2_MC1_v3_2[2]), .ZN(MCInst2_MC1_v3_3[0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[2]), .ZN(MCInst2_MC1_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_1_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        MCInst2_MC1_v0_3[0]), .Z(MCInst2_MC1_v0_0[1]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_1_U1 ( .A(MCInst2_MC1_v0_0[3]), .B(
        MCInst2_MC1_v0_3[3]), .Z(MCInst2_MC1_v0_1[1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U2 ( .A(MCInst2_MC1_v0_2Inst_1_n3), .B(
        MCInst2_MC1_v0_3[0]), .ZN(MCInst2_MC1_v0_2[1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_3[3]), .ZN(MCInst2_MC1_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_3[0]), .Z(MCInst2_MC1_v0_3[1]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_1_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        Red_MCInst2_MC1_v1_1_0_), .Z(MCInst2_MC1_v1_1[1]) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_1_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .Z(MCInst2_MC1_v1_2[1]) );
  XOR2_X1 MCInst2_MC1_v1_3Inst_1_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_0[3]), .Z(MCInst2_MC1_v1_3[1]) );
  XOR2_X1 MCInst2_MC1_v2_0Inst_1_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[0]), .Z(MCInst2_MC1_v2_0[1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U2 ( .A(MCInst2_MC1_v2_1Inst_1_n3), .B(
        MCInst2_MC1_v2_0[0]), .ZN(MCInst2_MC1_v2_1[1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U3 ( .A(MCInst2_MC1_v2_2Inst_1_n6), .B(
        MCInst2_MC1_v2_2Inst_1_n5), .ZN(MCInst2_MC1_v2_2[1]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        MCInst2_MC1_v2_0[0]), .ZN(MCInst2_MC1_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_1_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(MCInst2_MC1_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC1_v3_0Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_2[2]), .Z(MCInst2_MC1_v3_0[1]) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_1_0_), .Z(MCInst2_MC1_v3_1[1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U2 ( .A(MCInst2_MC1_v3_3Inst_1_n3), .B(
        MCInst2_MC1_v3_2[2]), .ZN(MCInst2_MC1_v3_3[1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_1_0_), .ZN(MCInst2_MC1_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_3[0]), .Z(MCInst2_MC1_v0_0[2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_2_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        MCInst2_MC1_v0_3[0]), .Z(MCInst2_MC1_v0_1[2]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_2_U1 ( .A(MCInst2_MC1_v0_0[3]), .B(
        MCInst2_MC1_v0_3[0]), .Z(MCInst2_MC1_v0_2[2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U2 ( .A(MCInst2_MC1_v1_1Inst_2_n3), .B(
        MCInst2_MC1_v1_0[3]), .ZN(MCInst2_MC1_v1_1[2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U2 ( .A(MCInst2_MC1_v1_2Inst_2_n3), .B(
        Red_MCInst2_MC1_v1_1_0_), .ZN(MCInst2_MC1_v1_2[2]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U2 ( .A(MCInst2_MC1_v2_1Inst_2_n3), .B(
        MCInst2_MC1_v2_0[0]), .ZN(MCInst2_MC1_v2_1[2]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U2 ( .A(MCInst2_MC1_v2_2Inst_2_n3), .B(
        MCInst2_MC1_v2_0[0]), .ZN(MCInst2_MC1_v2_2[2]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_2_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(MCInst2_MC1_v2_3[2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U2 ( .A(MCInst2_MC1_v3_1Inst_2_n3), .B(
        MCInst2_MC1_v3_2[2]), .ZN(MCInst2_MC1_v3_1[2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[2]), .ZN(MCInst2_MC1_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_2_U1 ( .A(MCInst2_MC1_v3_0[2]), .B(
        MCInst2_MC1_v3_2[2]), .Z(MCInst2_MC1_v3_3[2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_3[0]), .Z(MCInst2_MC1_v0_1[3]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_3[3]), .Z(MCInst2_MC1_v0_2[3]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_3_U1 ( .A(MCInst2_MC1_v1_3[2]), .B(
        Red_MCInst2_MC1_v1_1_0_), .Z(MCInst2_MC1_v1_1[3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U3 ( .A(MCInst2_MC1_v1_2Inst_3_n6), .B(
        MCInst2_MC1_v1_2Inst_3_n5), .ZN(MCInst2_MC1_v1_2[3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U2 ( .A(Red_MCInst2_MC1_v1_1_0_), .B(
        MCInst2_MC1_v1_0[3]), .ZN(MCInst2_MC1_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_3_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .Z(MCInst2_MC1_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_3_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[0]), .Z(MCInst2_MC1_v2_1[3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U2 ( .A(MCInst2_MC1_v2_2Inst_3_n3), .B(
        MCInst2_MC1_v2_0[0]), .ZN(MCInst2_MC1_v2_2[3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U2 ( .A(MCInst2_MC1_v2_3Inst_3_n3), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_3[3]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .ZN(MCInst2_MC1_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_3_U1 ( .A(MCInst2_MC1_v3_0[2]), .B(
        Red_MCInst2_MC1_v3_1_0_), .Z(MCInst2_MC1_v3_1[3]) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_3_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_1_0_), .Z(MCInst2_MC1_v3_3[3]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[56]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_0[0]), .B(
        MCInst2_MC1_v1_0[0]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        MCInst2_MC1_v3_2[2]), .Z(MCInst2_MC1_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[57]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_0[1]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_0[1]), .B(
        MCInst2_MC1_v3_0[1]), .Z(MCInst2_MC1_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[58]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_0[2]), .B(
        Red_MCInst2_MC1_v1_1_0_), .ZN(MCInst2_MC1_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_0[2]), .B(
        MCInst2_MC1_v3_0[2]), .Z(MCInst2_MC1_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[59]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        MCInst2_MC1_v1_0[3]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_0[3]), .B(
        Red_MCInst2_MC1_v3_1_0_), .Z(MCInst2_MC1_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[40]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_1[0]), .B(
        MCInst2_MC1_v1_1[0]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U1 ( .A(MCInst2_MC1_v0_0[3]), .B(
        MCInst2_MC1_v3_1[0]), .Z(MCInst2_MC1_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[41]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v1_1[1]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_1[1]), .B(
        MCInst2_MC1_v3_1[1]), .Z(MCInst2_MC1_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[42]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_1[2]), .B(
        MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_1[2]), .B(
        MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[43]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_1[3]), .B(
        MCInst2_MC1_v1_1[3]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_1[3]), .B(
        MCInst2_MC1_v3_1[3]), .Z(MCInst2_MC1_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[24]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_2[0]), .B(
        MCInst2_MC1_v1_2[0]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC1_v0_2[0]), .B(
        MCInst2_MC1_v3_2[0]), .Z(MCInst2_MC1_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[25]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_2[1]), .B(
        MCInst2_MC1_v1_2[1]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_2[1]), .B(
        Red_MCInst2_MC1_v3_1_0_), .Z(MCInst2_MC1_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[26]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_2[2]), .B(
        MCInst2_MC1_v1_2[2]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_2[2]), .B(
        MCInst2_MC1_v3_2[2]), .Z(MCInst2_MC1_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[27]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_2[3]), .B(
        MCInst2_MC1_v1_2[3]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_2[3]), .B(
        MCInst2_MC1_v3_2[3]), .Z(MCInst2_MC1_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[8]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_3[0]), .B(
        MCInst2_MC1_v1_0[3]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U1 ( .A(MCInst2_MC1_v0_3[0]), .B(
        MCInst2_MC1_v3_3[0]), .Z(MCInst2_MC1_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[9]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v1_3[1]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_3[1]), .B(
        MCInst2_MC1_v3_3[1]), .Z(MCInst2_MC1_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[10]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_3[2]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_0[3]), .B(
        MCInst2_MC1_v3_3[2]), .Z(MCInst2_MC1_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[11]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_3[3]), .B(
        Red_MCInst2_MC1_v1_1_0_), .ZN(MCInst2_MC1_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        MCInst2_MC1_v3_3[3]), .Z(MCInst2_MC1_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U2 ( .A(MCInst2_MC2_v0_2Inst_0_n3), .B(
        MCInst2_MC2_v0_3[0]), .ZN(MCInst2_MC2_v0_2[0]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_0[3]), .ZN(MCInst2_MC2_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_0_U1 ( .A(Red_MCInst2_MC2_v1_1_0_), .B(
        MCInst2_MC2_v1_0[3]), .Z(MCInst2_MC2_v1_1[0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U2 ( .A(MCInst2_MC2_v1_2Inst_0_n3), .B(
        MCInst2_MC2_v1_0[3]), .ZN(MCInst2_MC2_v1_2[0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U1 ( .A(MCInst2_MC2_v1_3[2]), .B(
        Red_MCInst2_MC2_v1_1_0_), .ZN(MCInst2_MC2_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_0_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[3]), .Z(MCInst2_MC2_v2_1[0]) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_0_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[0]), .Z(MCInst2_MC2_v2_2[0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U3 ( .A(MCInst2_MC2_v2_3Inst_0_n6), .B(
        MCInst2_MC2_v2_3Inst_0_n5), .ZN(MCInst2_MC2_v2_3[0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        MCInst2_MC2_v2_0[0]), .ZN(MCInst2_MC2_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_0_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(MCInst2_MC2_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_0_U1 ( .A(Red_MCInst2_MC2_v3_1_0_), .B(
        MCInst2_MC2_v3_2[2]), .Z(MCInst2_MC2_v3_1[0]) );
  XOR2_X1 MCInst2_MC2_v3_2Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[2]), .Z(MCInst2_MC2_v3_2[0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U2 ( .A(MCInst2_MC2_v3_3Inst_0_n3), .B(
        MCInst2_MC2_v3_2[2]), .ZN(MCInst2_MC2_v3_3[0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[2]), .ZN(MCInst2_MC2_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_1_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        MCInst2_MC2_v0_3[0]), .Z(MCInst2_MC2_v0_0[1]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_1_U1 ( .A(MCInst2_MC2_v0_0[3]), .B(
        MCInst2_MC2_v0_3[3]), .Z(MCInst2_MC2_v0_1[1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U2 ( .A(MCInst2_MC2_v0_2Inst_1_n3), .B(
        MCInst2_MC2_v0_3[0]), .ZN(MCInst2_MC2_v0_2[1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_3[3]), .ZN(MCInst2_MC2_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_3[0]), .Z(MCInst2_MC2_v0_3[1]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_1_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        Red_MCInst2_MC2_v1_1_0_), .Z(MCInst2_MC2_v1_1[1]) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_1_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .Z(MCInst2_MC2_v1_2[1]) );
  XOR2_X1 MCInst2_MC2_v1_3Inst_1_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_0[3]), .Z(MCInst2_MC2_v1_3[1]) );
  XOR2_X1 MCInst2_MC2_v2_0Inst_1_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[0]), .Z(MCInst2_MC2_v2_0[1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U2 ( .A(MCInst2_MC2_v2_1Inst_1_n3), .B(
        MCInst2_MC2_v2_0[0]), .ZN(MCInst2_MC2_v2_1[1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U3 ( .A(MCInst2_MC2_v2_2Inst_1_n6), .B(
        MCInst2_MC2_v2_2Inst_1_n5), .ZN(MCInst2_MC2_v2_2[1]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        MCInst2_MC2_v2_0[0]), .ZN(MCInst2_MC2_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_1_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(MCInst2_MC2_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC2_v3_0Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_2[2]), .Z(MCInst2_MC2_v3_0[1]) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_1_0_), .Z(MCInst2_MC2_v3_1[1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U2 ( .A(MCInst2_MC2_v3_3Inst_1_n3), .B(
        MCInst2_MC2_v3_2[2]), .ZN(MCInst2_MC2_v3_3[1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_1_0_), .ZN(MCInst2_MC2_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_3[0]), .Z(MCInst2_MC2_v0_0[2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_2_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        MCInst2_MC2_v0_3[0]), .Z(MCInst2_MC2_v0_1[2]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_2_U1 ( .A(MCInst2_MC2_v0_0[3]), .B(
        MCInst2_MC2_v0_3[0]), .Z(MCInst2_MC2_v0_2[2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U2 ( .A(MCInst2_MC2_v1_1Inst_2_n3), .B(
        MCInst2_MC2_v1_0[3]), .ZN(MCInst2_MC2_v1_1[2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U2 ( .A(MCInst2_MC2_v1_2Inst_2_n3), .B(
        Red_MCInst2_MC2_v1_1_0_), .ZN(MCInst2_MC2_v1_2[2]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U2 ( .A(MCInst2_MC2_v2_1Inst_2_n3), .B(
        MCInst2_MC2_v2_0[0]), .ZN(MCInst2_MC2_v2_1[2]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U2 ( .A(MCInst2_MC2_v2_2Inst_2_n3), .B(
        MCInst2_MC2_v2_0[0]), .ZN(MCInst2_MC2_v2_2[2]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_2_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(MCInst2_MC2_v2_3[2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U2 ( .A(MCInst2_MC2_v3_1Inst_2_n3), .B(
        MCInst2_MC2_v3_2[2]), .ZN(MCInst2_MC2_v3_1[2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[2]), .ZN(MCInst2_MC2_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_2_U1 ( .A(MCInst2_MC2_v3_0[2]), .B(
        MCInst2_MC2_v3_2[2]), .Z(MCInst2_MC2_v3_3[2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_3[0]), .Z(MCInst2_MC2_v0_1[3]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_3[3]), .Z(MCInst2_MC2_v0_2[3]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_3_U1 ( .A(MCInst2_MC2_v1_3[2]), .B(
        Red_MCInst2_MC2_v1_1_0_), .Z(MCInst2_MC2_v1_1[3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U3 ( .A(MCInst2_MC2_v1_2Inst_3_n6), .B(
        MCInst2_MC2_v1_2Inst_3_n5), .ZN(MCInst2_MC2_v1_2[3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U2 ( .A(Red_MCInst2_MC2_v1_1_0_), .B(
        MCInst2_MC2_v1_0[3]), .ZN(MCInst2_MC2_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_3_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .Z(MCInst2_MC2_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_3_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[0]), .Z(MCInst2_MC2_v2_1[3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U2 ( .A(MCInst2_MC2_v2_2Inst_3_n3), .B(
        MCInst2_MC2_v2_0[0]), .ZN(MCInst2_MC2_v2_2[3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U2 ( .A(MCInst2_MC2_v2_3Inst_3_n3), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_3[3]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .ZN(MCInst2_MC2_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_3_U1 ( .A(MCInst2_MC2_v3_0[2]), .B(
        Red_MCInst2_MC2_v3_1_0_), .Z(MCInst2_MC2_v3_1[3]) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_3_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_1_0_), .Z(MCInst2_MC2_v3_3[3]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[52]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_0[0]), .B(
        MCInst2_MC2_v1_0[0]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        MCInst2_MC2_v3_2[2]), .Z(MCInst2_MC2_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[53]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_0[1]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_0[1]), .B(
        MCInst2_MC2_v3_0[1]), .Z(MCInst2_MC2_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[54]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_0[2]), .B(
        Red_MCInst2_MC2_v1_1_0_), .ZN(MCInst2_MC2_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_0[2]), .B(
        MCInst2_MC2_v3_0[2]), .Z(MCInst2_MC2_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[55]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        MCInst2_MC2_v1_0[3]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_0[3]), .B(
        Red_MCInst2_MC2_v3_1_0_), .Z(MCInst2_MC2_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[36]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_1[0]), .B(
        MCInst2_MC2_v1_1[0]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U1 ( .A(MCInst2_MC2_v0_0[3]), .B(
        MCInst2_MC2_v3_1[0]), .Z(MCInst2_MC2_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[37]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v1_1[1]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_1[1]), .B(
        MCInst2_MC2_v3_1[1]), .Z(MCInst2_MC2_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[38]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_1[2]), .B(
        MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_1[2]), .B(
        MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[39]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_1[3]), .B(
        MCInst2_MC2_v1_1[3]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_1[3]), .B(
        MCInst2_MC2_v3_1[3]), .Z(MCInst2_MC2_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[20]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_2[0]), .B(
        MCInst2_MC2_v1_2[0]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC2_v0_2[0]), .B(
        MCInst2_MC2_v3_2[0]), .Z(MCInst2_MC2_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[21]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_2[1]), .B(
        MCInst2_MC2_v1_2[1]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_2[1]), .B(
        Red_MCInst2_MC2_v3_1_0_), .Z(MCInst2_MC2_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[22]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_2[2]), .B(
        MCInst2_MC2_v1_2[2]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_2[2]), .B(
        MCInst2_MC2_v3_2[2]), .Z(MCInst2_MC2_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[23]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_2[3]), .B(
        MCInst2_MC2_v1_2[3]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_2[3]), .B(
        MCInst2_MC2_v3_2[3]), .Z(MCInst2_MC2_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[4]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_3[0]), .B(
        MCInst2_MC2_v1_0[3]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U1 ( .A(MCInst2_MC2_v0_3[0]), .B(
        MCInst2_MC2_v3_3[0]), .Z(MCInst2_MC2_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[5]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v1_3[1]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_3[1]), .B(
        MCInst2_MC2_v3_3[1]), .Z(MCInst2_MC2_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[6]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_3[2]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_0[3]), .B(
        MCInst2_MC2_v3_3[2]), .Z(MCInst2_MC2_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[7]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_3[3]), .B(
        Red_MCInst2_MC2_v1_1_0_), .ZN(MCInst2_MC2_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        MCInst2_MC2_v3_3[3]), .Z(MCInst2_MC2_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U2 ( .A(MCInst2_MC3_v0_2Inst_0_n3), .B(
        MCInst2_MC3_v0_3[0]), .ZN(MCInst2_MC3_v0_2[0]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_0[3]), .ZN(MCInst2_MC3_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_0_U1 ( .A(Red_MCInst2_MC3_v1_1_0_), .B(
        MCInst2_MC3_v1_0[3]), .Z(MCInst2_MC3_v1_1[0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U2 ( .A(MCInst2_MC3_v1_2Inst_0_n3), .B(
        MCInst2_MC3_v1_0[3]), .ZN(MCInst2_MC3_v1_2[0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U1 ( .A(MCInst2_MC3_v1_3[2]), .B(
        Red_MCInst2_MC3_v1_1_0_), .ZN(MCInst2_MC3_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_0_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[3]), .Z(MCInst2_MC3_v2_1[0]) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_0_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[0]), .Z(MCInst2_MC3_v2_2[0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U3 ( .A(MCInst2_MC3_v2_3Inst_0_n6), .B(
        MCInst2_MC3_v2_3Inst_0_n5), .ZN(MCInst2_MC3_v2_3[0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        MCInst2_MC3_v2_0[0]), .ZN(MCInst2_MC3_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_0_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(MCInst2_MC3_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_0_U1 ( .A(Red_MCInst2_MC3_v3_1_0_), .B(
        MCInst2_MC3_v3_2[2]), .Z(MCInst2_MC3_v3_1[0]) );
  XOR2_X1 MCInst2_MC3_v3_2Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[2]), .Z(MCInst2_MC3_v3_2[0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U2 ( .A(MCInst2_MC3_v3_3Inst_0_n3), .B(
        MCInst2_MC3_v3_2[2]), .ZN(MCInst2_MC3_v3_3[0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[2]), .ZN(MCInst2_MC3_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_1_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        MCInst2_MC3_v0_3[0]), .Z(MCInst2_MC3_v0_0[1]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_1_U1 ( .A(MCInst2_MC3_v0_0[3]), .B(
        MCInst2_MC3_v0_3[3]), .Z(MCInst2_MC3_v0_1[1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U2 ( .A(MCInst2_MC3_v0_2Inst_1_n3), .B(
        MCInst2_MC3_v0_3[0]), .ZN(MCInst2_MC3_v0_2[1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_3[3]), .ZN(MCInst2_MC3_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_3[0]), .Z(MCInst2_MC3_v0_3[1]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_1_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        Red_MCInst2_MC3_v1_1_0_), .Z(MCInst2_MC3_v1_1[1]) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_1_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .Z(MCInst2_MC3_v1_2[1]) );
  XOR2_X1 MCInst2_MC3_v1_3Inst_1_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_0[3]), .Z(MCInst2_MC3_v1_3[1]) );
  XOR2_X1 MCInst2_MC3_v2_0Inst_1_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[0]), .Z(MCInst2_MC3_v2_0[1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U2 ( .A(MCInst2_MC3_v2_1Inst_1_n3), .B(
        MCInst2_MC3_v2_0[0]), .ZN(MCInst2_MC3_v2_1[1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U3 ( .A(MCInst2_MC3_v2_2Inst_1_n6), .B(
        MCInst2_MC3_v2_2Inst_1_n5), .ZN(MCInst2_MC3_v2_2[1]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        MCInst2_MC3_v2_0[0]), .ZN(MCInst2_MC3_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_1_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(MCInst2_MC3_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC3_v3_0Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_2[2]), .Z(MCInst2_MC3_v3_0[1]) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_1_0_), .Z(MCInst2_MC3_v3_1[1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U2 ( .A(MCInst2_MC3_v3_3Inst_1_n3), .B(
        MCInst2_MC3_v3_2[2]), .ZN(MCInst2_MC3_v3_3[1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_1_0_), .ZN(MCInst2_MC3_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_3[0]), .Z(MCInst2_MC3_v0_0[2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_2_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        MCInst2_MC3_v0_3[0]), .Z(MCInst2_MC3_v0_1[2]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_2_U1 ( .A(MCInst2_MC3_v0_0[3]), .B(
        MCInst2_MC3_v0_3[0]), .Z(MCInst2_MC3_v0_2[2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U2 ( .A(MCInst2_MC3_v1_1Inst_2_n3), .B(
        MCInst2_MC3_v1_0[3]), .ZN(MCInst2_MC3_v1_1[2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U2 ( .A(MCInst2_MC3_v1_2Inst_2_n3), .B(
        Red_MCInst2_MC3_v1_1_0_), .ZN(MCInst2_MC3_v1_2[2]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U2 ( .A(MCInst2_MC3_v2_1Inst_2_n3), .B(
        MCInst2_MC3_v2_0[0]), .ZN(MCInst2_MC3_v2_1[2]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U2 ( .A(MCInst2_MC3_v2_2Inst_2_n3), .B(
        MCInst2_MC3_v2_0[0]), .ZN(MCInst2_MC3_v2_2[2]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_2_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(MCInst2_MC3_v2_3[2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U2 ( .A(MCInst2_MC3_v3_1Inst_2_n3), .B(
        MCInst2_MC3_v3_2[2]), .ZN(MCInst2_MC3_v3_1[2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[2]), .ZN(MCInst2_MC3_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_2_U1 ( .A(MCInst2_MC3_v3_0[2]), .B(
        MCInst2_MC3_v3_2[2]), .Z(MCInst2_MC3_v3_3[2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_3[0]), .Z(MCInst2_MC3_v0_1[3]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_3[3]), .Z(MCInst2_MC3_v0_2[3]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_3_U1 ( .A(MCInst2_MC3_v1_3[2]), .B(
        Red_MCInst2_MC3_v1_1_0_), .Z(MCInst2_MC3_v1_1[3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U3 ( .A(MCInst2_MC3_v1_2Inst_3_n6), .B(
        MCInst2_MC3_v1_2Inst_3_n5), .ZN(MCInst2_MC3_v1_2[3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U2 ( .A(Red_MCInst2_MC3_v1_1_0_), .B(
        MCInst2_MC3_v1_0[3]), .ZN(MCInst2_MC3_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_3_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .Z(MCInst2_MC3_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_3_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[0]), .Z(MCInst2_MC3_v2_1[3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U2 ( .A(MCInst2_MC3_v2_2Inst_3_n3), .B(
        MCInst2_MC3_v2_0[0]), .ZN(MCInst2_MC3_v2_2[3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U2 ( .A(MCInst2_MC3_v2_3Inst_3_n3), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_3[3]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .ZN(MCInst2_MC3_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_3_U1 ( .A(MCInst2_MC3_v3_0[2]), .B(
        Red_MCInst2_MC3_v3_1_0_), .Z(MCInst2_MC3_v3_1[3]) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_3_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_1_0_), .Z(MCInst2_MC3_v3_3[3]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[48]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_0[0]), .B(
        MCInst2_MC3_v1_0[0]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        MCInst2_MC3_v3_2[2]), .Z(MCInst2_MC3_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[49]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_0[1]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_0[1]), .B(
        MCInst2_MC3_v3_0[1]), .Z(MCInst2_MC3_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[50]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_0[2]), .B(
        Red_MCInst2_MC3_v1_1_0_), .ZN(MCInst2_MC3_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_0[2]), .B(
        MCInst2_MC3_v3_0[2]), .Z(MCInst2_MC3_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[51]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        MCInst2_MC3_v1_0[3]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_0[3]), .B(
        Red_MCInst2_MC3_v3_1_0_), .Z(MCInst2_MC3_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[32]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_1[0]), .B(
        MCInst2_MC3_v1_1[0]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U1 ( .A(MCInst2_MC3_v0_0[3]), .B(
        MCInst2_MC3_v3_1[0]), .Z(MCInst2_MC3_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[33]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v1_1[1]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_1[1]), .B(
        MCInst2_MC3_v3_1[1]), .Z(MCInst2_MC3_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[34]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_1[2]), .B(
        MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_1[2]), .B(
        MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[35]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_1[3]), .B(
        MCInst2_MC3_v1_1[3]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_1[3]), .B(
        MCInst2_MC3_v3_1[3]), .Z(MCInst2_MC3_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[16]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_2[0]), .B(
        MCInst2_MC3_v1_2[0]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC3_v0_2[0]), .B(
        MCInst2_MC3_v3_2[0]), .Z(MCInst2_MC3_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[17]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_2[1]), .B(
        MCInst2_MC3_v1_2[1]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_2[1]), .B(
        Red_MCInst2_MC3_v3_1_0_), .Z(MCInst2_MC3_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[18]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_2[2]), .B(
        MCInst2_MC3_v1_2[2]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_2[2]), .B(
        MCInst2_MC3_v3_2[2]), .Z(MCInst2_MC3_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[19]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_2[3]), .B(
        MCInst2_MC3_v1_2[3]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_2[3]), .B(
        MCInst2_MC3_v3_2[3]), .Z(MCInst2_MC3_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[0]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_3[0]), .B(
        MCInst2_MC3_v1_0[3]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U1 ( .A(MCInst2_MC3_v0_3[0]), .B(
        MCInst2_MC3_v3_3[0]), .Z(MCInst2_MC3_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[1]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v1_3[1]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_3[1]), .B(
        MCInst2_MC3_v3_3[1]), .Z(MCInst2_MC3_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[2]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_3[2]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_0[3]), .B(
        MCInst2_MC3_v3_3[2]), .Z(MCInst2_MC3_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[3]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_3[3]), .B(
        Red_MCInst2_MC3_v1_1_0_), .ZN(MCInst2_MC3_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        MCInst2_MC3_v3_3[3]), .Z(MCInst2_MC3_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_0_LFInst_0_n5), .ZN(Red_Plaintext[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(Plaintext[2]), .B(
        Plaintext[3]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Plaintext[0]), .B(
        Plaintext[1]), .Z(Red_PlaintextInst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_1_LFInst_0_n5), .ZN(Red_Plaintext[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(Plaintext[6]), .B(
        Plaintext[7]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Plaintext[4]), .B(
        Plaintext[5]), .Z(Red_PlaintextInst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_2_LFInst_0_n5), .ZN(Red_Plaintext[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(Plaintext[10]), .B(
        Plaintext[11]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Plaintext[8]), .B(
        Plaintext[9]), .Z(Red_PlaintextInst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_3_LFInst_0_n5), .ZN(Red_Plaintext[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(Plaintext[14]), .B(
        Plaintext[15]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Plaintext[12]), .B(
        Plaintext[13]), .Z(Red_PlaintextInst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_4_LFInst_0_n5), .ZN(Red_Plaintext[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(Plaintext[18]), .B(
        Plaintext[19]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Plaintext[16]), .B(
        Plaintext[17]), .Z(Red_PlaintextInst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_5_LFInst_0_n5), .ZN(Red_Plaintext[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(Plaintext[22]), .B(
        Plaintext[23]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Plaintext[20]), .B(
        Plaintext[21]), .Z(Red_PlaintextInst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_6_LFInst_0_n5), .ZN(Red_Plaintext[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(Plaintext[26]), .B(
        Plaintext[27]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Plaintext[24]), .B(
        Plaintext[25]), .Z(Red_PlaintextInst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_7_LFInst_0_n5), .ZN(Red_Plaintext[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(Plaintext[30]), .B(
        Plaintext[31]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Plaintext[28]), .B(
        Plaintext[29]), .Z(Red_PlaintextInst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_8_LFInst_0_n5), .ZN(Red_Plaintext[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(Plaintext[34]), .B(
        Plaintext[35]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Plaintext[32]), .B(
        Plaintext[33]), .Z(Red_PlaintextInst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_9_LFInst_0_n5), .ZN(Red_Plaintext[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(Plaintext[38]), .B(
        Plaintext[39]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Plaintext[36]), .B(
        Plaintext[37]), .Z(Red_PlaintextInst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_10_LFInst_0_n5), .ZN(Red_Plaintext[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(Plaintext[42]), .B(
        Plaintext[43]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Plaintext[40]), .B(
        Plaintext[41]), .Z(Red_PlaintextInst_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_11_LFInst_0_n5), .ZN(Red_Plaintext[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(Plaintext[46]), .B(
        Plaintext[47]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Plaintext[44]), .B(
        Plaintext[45]), .Z(Red_PlaintextInst_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_12_LFInst_0_n5), .ZN(Red_Plaintext[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(Plaintext[50]), .B(
        Plaintext[51]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Plaintext[48]), .B(
        Plaintext[49]), .Z(Red_PlaintextInst_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_13_LFInst_0_n5), .ZN(Red_Plaintext[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(Plaintext[54]), .B(
        Plaintext[55]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Plaintext[52]), .B(
        Plaintext[53]), .Z(Red_PlaintextInst_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_14_LFInst_0_n5), .ZN(Red_Plaintext[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(Plaintext[58]), .B(
        Plaintext[59]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Plaintext[56]), .B(
        Plaintext[57]), .Z(Red_PlaintextInst_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_15_LFInst_0_n5), .ZN(Red_Plaintext[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(Plaintext[62]), .B(
        Plaintext[63]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Plaintext[60]), .B(
        Plaintext[61]), .Z(Red_PlaintextInst_LFInst_15_LFInst_0_n6) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_0_U1 ( .A(Red_Plaintext[0]), .B(
        Red_RoundKey[0]), .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_0_U1 ( .A(Red_Plaintext[1]), .B(
        Red_RoundKey[1]), .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_0_U1 ( .A(Red_Plaintext[2]), .B(
        Red_RoundKey[2]), .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_0_U1 ( .A(Red_Plaintext[3]), .B(
        Red_RoundKey[3]), .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_0_U1 ( .A(Red_Plaintext[4]), .B(
        Red_RoundKey[4]), .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_0_U1 ( .A(Red_Plaintext[5]), .B(
        Red_RoundKey[5]), .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_0_U1 ( .A(Red_Plaintext[6]), .B(
        Red_RoundKey[6]), .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_0_U1 ( .A(Red_Plaintext[7]), .B(
        Red_RoundKey[7]), .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_0_U1 ( .A(Red_Plaintext[8]), .B(
        Red_RoundKey[8]), .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_0_U1 ( .A(Red_Plaintext[9]), .B(
        Red_RoundKey[9]), .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_0_U1 ( .A(Red_Plaintext[10]), .B(
        Red_RoundKey[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_0_U1 ( .A(Red_Plaintext[11]), .B(
        Red_RoundKey[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_0_U1 ( .A(Red_Plaintext[12]), .B(
        Red_RoundKey[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_0_U1 ( .A(Red_Plaintext[13]), .B(
        Red_RoundKey[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_0_U1 ( .A(Red_Plaintext[14]), .B(
        Red_RoundKey[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_0_U1 ( .A(Red_Plaintext[15]), .B(
        Red_RoundKey[15]), .Z(Red_AddRoundKeyOutput[15]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[3]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U3 ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U2 ( .A1(AddRoundKeyOutput[3]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U1 ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[0]) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U3 ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U2 ( .A1(AddRoundKeyOutput[7]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U1 ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[1]) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U3 ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U2 ( .A1(AddRoundKeyOutput[11]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U1 ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[2]) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U3 ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U2 ( .A1(AddRoundKeyOutput[15]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U1 ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_4_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[6]) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U2 ( .A1(AddRoundKeyOutput[19]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U1 ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_5_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[7]) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U2 ( .A1(AddRoundKeyOutput[23]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U1 ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_6_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[4]) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U2 ( .A1(AddRoundKeyOutput[27]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U1 ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_7_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[5]) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U2 ( .A1(AddRoundKeyOutput[31]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U1 ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[9]) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U3 ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U2 ( .A1(AddRoundKeyOutput[35]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U1 ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[10]) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U3 ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U2 ( .A1(AddRoundKeyOutput[39]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U1 ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[11])
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U3 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U2 ( .A1(AddRoundKeyOutput[43]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U1 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[8]) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U3 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U2 ( .A1(AddRoundKeyOutput[47]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U1 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[12])
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U3 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U2 ( .A1(AddRoundKeyOutput[51]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U1 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[13])
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U2 ( .A1(AddRoundKeyOutput[55]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U1 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[14])
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U3 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U2 ( .A1(AddRoundKeyOutput[59]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U1 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n7)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n9), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n8), .ZN(Red_ShiftRowsOutput[15])
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U3 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n8)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U2 ( .A1(AddRoundKeyOutput[63]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_0_n7), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U1 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_v0_0Inst_0_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_0[3]), .Z(Red_MCInst_MC0_v0_0_0_) );
  XOR2_X1 Red_MCInst_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_3[0]), .Z(Red_MCInst_MC0_v0_2_0_) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_0_U2 ( .A(Red_MCInst_MC0_v0_3Inst_0_n3), 
        .B(MCInst_MC0_v0_3[3]), .ZN(Red_MCInst_MC0_v0_3_0_) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_0_U1 ( .A(Red_MCInst_MC0_v0_1_0_), .B(
        MCInst_MC0_v0_0[3]), .ZN(Red_MCInst_MC0_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U3 ( .A(Red_MCInst_MC0_v1_0Inst_0_n6), 
        .B(Red_MCInst_MC0_v1_0Inst_0_n5), .ZN(Red_MCInst_MC0_v1_0_0_) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U2 ( .A(Red_MCInst_MC0_v1_1_0_), .B(
        MCInst_MC0_v1_0[3]), .ZN(Red_MCInst_MC0_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .Z(Red_MCInst_MC0_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC0_v1_2Inst_0_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        Red_MCInst_MC0_v1_1_0_), .Z(Red_MCInst_MC0_v1_2_0_) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_0_U2 ( .A(Red_MCInst_MC0_v1_3Inst_0_n3), 
        .B(Red_MCInst_MC0_v1_1_0_), .ZN(Red_MCInst_MC0_v1_3_0_) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_0_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .ZN(Red_MCInst_MC0_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_0_U2 ( .A(Red_MCInst_MC0_v2_0Inst_0_n3), 
        .B(MCInst_MC0_v2_0[3]), .ZN(Red_MCInst_MC0_v2_0_0_) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .ZN(Red_MCInst_MC0_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC0_v2_1Inst_0_U1 ( .A(MCInst_MC0_v2_0[3]), .B(
        MCInst_MC0_v2_0[0]), .Z(Red_MCInst_MC0_v2_1_0_) );
  XOR2_X1 Red_MCInst_MC0_v2_2Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_2_0_) );
  XOR2_X1 Red_MCInst_MC0_v2_3Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[0]), .Z(Red_MCInst_MC0_v2_3_0_) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_0_U2 ( .A(Red_MCInst_MC0_v3_0Inst_0_n3), 
        .B(Red_MCInst_MC0_v3_1_0_), .ZN(Red_MCInst_MC0_v3_0_0_) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[2]), .ZN(Red_MCInst_MC0_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U2 ( .A(Red_MCInst_MC0_v3_2Inst_0_n3), 
        .B(MCInst_MC0_v3_2[2]), .ZN(Red_MCInst_MC0_v3_2_0_) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U1 ( .A(MCInst_MC0_v3_0[2]), .B(
        Red_MCInst_MC0_v3_1_0_), .ZN(Red_MCInst_MC0_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC0_v3_3Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_2[2]), .Z(Red_MCInst_MC0_v3_3_0_) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[15]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_0_0_), 
        .B(Red_MCInst_MC0_v1_0_0_), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_0_0_), 
        .B(Red_MCInst_MC0_v3_0_0_), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[11]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_1_0_), 
        .B(Red_MCInst_MC0_v1_1_0_), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_1_0_), 
        .B(Red_MCInst_MC0_v3_1_0_), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[7]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_2_0_), 
        .B(Red_MCInst_MC0_v1_2_0_), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_2_0_), 
        .B(Red_MCInst_MC0_v3_2_0_), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[3]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_3_0_), 
        .B(Red_MCInst_MC0_v1_3_0_), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_3_0_), 
        .B(Red_MCInst_MC0_v3_3_0_), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_0_n8)
         );
  XOR2_X1 Red_MCInst_MC1_v0_0Inst_0_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_0[3]), .Z(Red_MCInst_MC1_v0_0_0_) );
  XOR2_X1 Red_MCInst_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_3[0]), .Z(Red_MCInst_MC1_v0_2_0_) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_0_U2 ( .A(Red_MCInst_MC1_v0_3Inst_0_n3), 
        .B(MCInst_MC1_v0_3[3]), .ZN(Red_MCInst_MC1_v0_3_0_) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_0_U1 ( .A(Red_MCInst_MC1_v0_1_0_), .B(
        MCInst_MC1_v0_0[3]), .ZN(Red_MCInst_MC1_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U3 ( .A(Red_MCInst_MC1_v1_0Inst_0_n6), 
        .B(Red_MCInst_MC1_v1_0Inst_0_n5), .ZN(Red_MCInst_MC1_v1_0_0_) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U2 ( .A(Red_MCInst_MC1_v1_1_0_), .B(
        MCInst_MC1_v1_0[3]), .ZN(Red_MCInst_MC1_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .Z(Red_MCInst_MC1_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC1_v1_2Inst_0_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        Red_MCInst_MC1_v1_1_0_), .Z(Red_MCInst_MC1_v1_2_0_) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_0_U2 ( .A(Red_MCInst_MC1_v1_3Inst_0_n3), 
        .B(Red_MCInst_MC1_v1_1_0_), .ZN(Red_MCInst_MC1_v1_3_0_) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_0_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .ZN(Red_MCInst_MC1_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_0_U2 ( .A(Red_MCInst_MC1_v2_0Inst_0_n3), 
        .B(MCInst_MC1_v2_0[3]), .ZN(Red_MCInst_MC1_v2_0_0_) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .ZN(Red_MCInst_MC1_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC1_v2_1Inst_0_U1 ( .A(MCInst_MC1_v2_0[3]), .B(
        MCInst_MC1_v2_0[0]), .Z(Red_MCInst_MC1_v2_1_0_) );
  XOR2_X1 Red_MCInst_MC1_v2_2Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_2_0_) );
  XOR2_X1 Red_MCInst_MC1_v2_3Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[0]), .Z(Red_MCInst_MC1_v2_3_0_) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_0_U2 ( .A(Red_MCInst_MC1_v3_0Inst_0_n3), 
        .B(Red_MCInst_MC1_v3_1_0_), .ZN(Red_MCInst_MC1_v3_0_0_) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[2]), .ZN(Red_MCInst_MC1_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U2 ( .A(Red_MCInst_MC1_v3_2Inst_0_n3), 
        .B(MCInst_MC1_v3_2[2]), .ZN(Red_MCInst_MC1_v3_2_0_) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U1 ( .A(MCInst_MC1_v3_0[2]), .B(
        Red_MCInst_MC1_v3_1_0_), .ZN(Red_MCInst_MC1_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC1_v3_3Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_2[2]), .Z(Red_MCInst_MC1_v3_3_0_) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[14]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_0_0_), 
        .B(Red_MCInst_MC1_v1_0_0_), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_0_0_), 
        .B(Red_MCInst_MC1_v3_0_0_), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[10]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_1_0_), 
        .B(Red_MCInst_MC1_v1_1_0_), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_1_0_), 
        .B(Red_MCInst_MC1_v3_1_0_), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[6]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_2_0_), 
        .B(Red_MCInst_MC1_v1_2_0_), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_2_0_), 
        .B(Red_MCInst_MC1_v3_2_0_), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[2]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_3_0_), 
        .B(Red_MCInst_MC1_v1_3_0_), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_3_0_), 
        .B(Red_MCInst_MC1_v3_3_0_), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_0_n8)
         );
  XOR2_X1 Red_MCInst_MC2_v0_0Inst_0_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_0[3]), .Z(Red_MCInst_MC2_v0_0_0_) );
  XOR2_X1 Red_MCInst_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_3[0]), .Z(Red_MCInst_MC2_v0_2_0_) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_0_U2 ( .A(Red_MCInst_MC2_v0_3Inst_0_n3), 
        .B(MCInst_MC2_v0_3[3]), .ZN(Red_MCInst_MC2_v0_3_0_) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_0_U1 ( .A(Red_MCInst_MC2_v0_1_0_), .B(
        MCInst_MC2_v0_0[3]), .ZN(Red_MCInst_MC2_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U3 ( .A(Red_MCInst_MC2_v1_0Inst_0_n6), 
        .B(Red_MCInst_MC2_v1_0Inst_0_n5), .ZN(Red_MCInst_MC2_v1_0_0_) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U2 ( .A(Red_MCInst_MC2_v1_1_0_), .B(
        MCInst_MC2_v1_0[3]), .ZN(Red_MCInst_MC2_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .Z(Red_MCInst_MC2_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC2_v1_2Inst_0_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        Red_MCInst_MC2_v1_1_0_), .Z(Red_MCInst_MC2_v1_2_0_) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_0_U2 ( .A(Red_MCInst_MC2_v1_3Inst_0_n3), 
        .B(Red_MCInst_MC2_v1_1_0_), .ZN(Red_MCInst_MC2_v1_3_0_) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_0_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .ZN(Red_MCInst_MC2_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_0_U2 ( .A(Red_MCInst_MC2_v2_0Inst_0_n3), 
        .B(MCInst_MC2_v2_0[3]), .ZN(Red_MCInst_MC2_v2_0_0_) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .ZN(Red_MCInst_MC2_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC2_v2_1Inst_0_U1 ( .A(MCInst_MC2_v2_0[3]), .B(
        MCInst_MC2_v2_0[0]), .Z(Red_MCInst_MC2_v2_1_0_) );
  XOR2_X1 Red_MCInst_MC2_v2_2Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_2_0_) );
  XOR2_X1 Red_MCInst_MC2_v2_3Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[0]), .Z(Red_MCInst_MC2_v2_3_0_) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_0_U2 ( .A(Red_MCInst_MC2_v3_0Inst_0_n3), 
        .B(Red_MCInst_MC2_v3_1_0_), .ZN(Red_MCInst_MC2_v3_0_0_) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[2]), .ZN(Red_MCInst_MC2_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U2 ( .A(Red_MCInst_MC2_v3_2Inst_0_n3), 
        .B(MCInst_MC2_v3_2[2]), .ZN(Red_MCInst_MC2_v3_2_0_) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U1 ( .A(MCInst_MC2_v3_0[2]), .B(
        Red_MCInst_MC2_v3_1_0_), .ZN(Red_MCInst_MC2_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC2_v3_3Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_2[2]), .Z(Red_MCInst_MC2_v3_3_0_) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[13]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_0_0_), 
        .B(Red_MCInst_MC2_v1_0_0_), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_0_0_), 
        .B(Red_MCInst_MC2_v3_0_0_), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[9]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_1_0_), 
        .B(Red_MCInst_MC2_v1_1_0_), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_1_0_), 
        .B(Red_MCInst_MC2_v3_1_0_), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[5]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_2_0_), 
        .B(Red_MCInst_MC2_v1_2_0_), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_2_0_), 
        .B(Red_MCInst_MC2_v3_2_0_), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[1]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_3_0_), 
        .B(Red_MCInst_MC2_v1_3_0_), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_3_0_), 
        .B(Red_MCInst_MC2_v3_3_0_), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_0_n8)
         );
  XOR2_X1 Red_MCInst_MC3_v0_0Inst_0_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_0[3]), .Z(Red_MCInst_MC3_v0_0_0_) );
  XOR2_X1 Red_MCInst_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_3[0]), .Z(Red_MCInst_MC3_v0_2_0_) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_0_U2 ( .A(Red_MCInst_MC3_v0_3Inst_0_n3), 
        .B(MCInst_MC3_v0_3[3]), .ZN(Red_MCInst_MC3_v0_3_0_) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_0_U1 ( .A(Red_MCInst_MC3_v0_1_0_), .B(
        MCInst_MC3_v0_0[3]), .ZN(Red_MCInst_MC3_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U3 ( .A(Red_MCInst_MC3_v1_0Inst_0_n6), 
        .B(Red_MCInst_MC3_v1_0Inst_0_n5), .ZN(Red_MCInst_MC3_v1_0_0_) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U2 ( .A(Red_MCInst_MC3_v1_1_0_), .B(
        MCInst_MC3_v1_0[3]), .ZN(Red_MCInst_MC3_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .Z(Red_MCInst_MC3_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC3_v1_2Inst_0_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        Red_MCInst_MC3_v1_1_0_), .Z(Red_MCInst_MC3_v1_2_0_) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_0_U2 ( .A(Red_MCInst_MC3_v1_3Inst_0_n3), 
        .B(Red_MCInst_MC3_v1_1_0_), .ZN(Red_MCInst_MC3_v1_3_0_) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_0_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .ZN(Red_MCInst_MC3_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_0_U2 ( .A(Red_MCInst_MC3_v2_0Inst_0_n3), 
        .B(MCInst_MC3_v2_0[3]), .ZN(Red_MCInst_MC3_v2_0_0_) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .ZN(Red_MCInst_MC3_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC3_v2_1Inst_0_U1 ( .A(MCInst_MC3_v2_0[3]), .B(
        MCInst_MC3_v2_0[0]), .Z(Red_MCInst_MC3_v2_1_0_) );
  XOR2_X1 Red_MCInst_MC3_v2_2Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_2_0_) );
  XOR2_X1 Red_MCInst_MC3_v2_3Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[0]), .Z(Red_MCInst_MC3_v2_3_0_) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_0_U2 ( .A(Red_MCInst_MC3_v3_0Inst_0_n3), 
        .B(Red_MCInst_MC3_v3_1_0_), .ZN(Red_MCInst_MC3_v3_0_0_) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[2]), .ZN(Red_MCInst_MC3_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U2 ( .A(Red_MCInst_MC3_v3_2Inst_0_n3), 
        .B(MCInst_MC3_v3_2[2]), .ZN(Red_MCInst_MC3_v3_2_0_) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U1 ( .A(MCInst_MC3_v3_0[2]), .B(
        Red_MCInst_MC3_v3_1_0_), .ZN(Red_MCInst_MC3_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC3_v3_3Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_2[2]), .Z(Red_MCInst_MC3_v3_3_0_) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[12]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_0_0_), 
        .B(Red_MCInst_MC3_v1_0_0_), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_0_0_), 
        .B(Red_MCInst_MC3_v3_0_0_), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[8]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_1_0_), 
        .B(Red_MCInst_MC3_v1_1_0_), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_1_0_), 
        .B(Red_MCInst_MC3_v3_1_0_), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[4]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_2_0_), 
        .B(Red_MCInst_MC3_v1_2_0_), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_2_0_), 
        .B(Red_MCInst_MC3_v3_2_0_), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[0]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_3_0_), 
        .B(Red_MCInst_MC3_v1_3_0_), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_3_0_), 
        .B(Red_MCInst_MC3_v3_3_0_), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_0_n8)
         );
  DFF_X1 RedStateReg_s_current_state_reg_0_ ( .D(Red_MC_output[0]), .CK(clk), 
        .Q(Red_SubCellInput2[0]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_1_ ( .D(Red_MC_output[1]), .CK(clk), 
        .Q(Red_SubCellInput2[1]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_2_ ( .D(Red_MC_output[2]), .CK(clk), 
        .Q(Red_SubCellInput2[2]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_3_ ( .D(Red_MC_output[3]), .CK(clk), 
        .Q(Red_SubCellInput2[3]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_4_ ( .D(Red_MC_output[4]), .CK(clk), 
        .Q(Red_SubCellInput2[4]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_5_ ( .D(Red_MC_output[5]), .CK(clk), 
        .Q(Red_SubCellInput2[5]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_6_ ( .D(Red_MC_output[6]), .CK(clk), 
        .Q(Red_SubCellInput2[6]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_7_ ( .D(Red_MC_output[7]), .CK(clk), 
        .Q(Red_SubCellInput2[7]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_8_ ( .D(Red_MC_output[8]), .CK(clk), 
        .Q(Red_SubCellInput2[8]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_9_ ( .D(Red_MC_output[9]), .CK(clk), 
        .Q(Red_SubCellInput2[9]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_10_ ( .D(Red_MC_output[10]), .CK(clk), 
        .Q(Red_SubCellInput2[10]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_11_ ( .D(Red_MC_output[11]), .CK(clk), 
        .Q(Red_SubCellInput2[11]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_12_ ( .D(Red_MC_output[12]), .CK(clk), 
        .Q(Red_SubCellInput2[12]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_13_ ( .D(Red_MC_output[13]), .CK(clk), 
        .Q(Red_SubCellInput2[13]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_14_ ( .D(Red_MC_output[14]), .CK(clk), 
        .Q(Red_SubCellInput2[14]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_15_ ( .D(Red_MC_output[15]), .CK(clk), 
        .Q(Red_SubCellInput2[15]), .QN() );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[3])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U3 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U2 ( .A1(SubCellInput2[3]), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U1 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[0])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U3 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U2 ( .A1(SubCellInput2[7]), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U1 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[1])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U3 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U2 ( .A1(SubCellInput2[11]), 
        .A2(Red_SubCellInst2_LFInst_2_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U1 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[2])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U3 ( .A1(SubCellInput2[12]), 
        .A2(SubCellInput2[13]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U2 ( .A1(SubCellInput2[15]), 
        .A2(Red_SubCellInst2_LFInst_3_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U1 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[6])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U3 ( .A1(SubCellInput2[16]), 
        .A2(SubCellInput2[17]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U2 ( .A1(SubCellInput2[19]), 
        .A2(Red_SubCellInst2_LFInst_4_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U1 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[18]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[7])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U3 ( .A1(SubCellInput2[20]), 
        .A2(SubCellInput2[21]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U2 ( .A1(SubCellInput2[23]), 
        .A2(Red_SubCellInst2_LFInst_5_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U1 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[22]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[4])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U3 ( .A1(SubCellInput2[24]), 
        .A2(SubCellInput2[25]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U2 ( .A1(SubCellInput2[27]), 
        .A2(Red_SubCellInst2_LFInst_6_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U1 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[26]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[5])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U3 ( .A1(SubCellInput2[28]), 
        .A2(SubCellInput2[29]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U2 ( .A1(SubCellInput2[31]), 
        .A2(Red_SubCellInst2_LFInst_7_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U1 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[30]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[9])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U3 ( .A1(SubCellInput2[32]), 
        .A2(SubCellInput2[33]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U2 ( .A1(SubCellInput2[35]), 
        .A2(Red_SubCellInst2_LFInst_8_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U1 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[34]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[10])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U3 ( .A1(SubCellInput2[36]), 
        .A2(SubCellInput2[37]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U2 ( .A1(SubCellInput2[39]), 
        .A2(Red_SubCellInst2_LFInst_9_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U1 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[38]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[11])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U3 ( .A1(SubCellInput2[40]), 
        .A2(SubCellInput2[41]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U2 ( .A1(SubCellInput2[43]), 
        .A2(Red_SubCellInst2_LFInst_10_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U1 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[42]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[8])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U3 ( .A1(SubCellInput2[44]), 
        .A2(SubCellInput2[45]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U2 ( .A1(SubCellInput2[47]), 
        .A2(Red_SubCellInst2_LFInst_11_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U1 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[12])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U3 ( .A1(SubCellInput2[48]), 
        .A2(SubCellInput2[49]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U2 ( .A1(SubCellInput2[51]), 
        .A2(Red_SubCellInst2_LFInst_12_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U1 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[50]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[13])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U3 ( .A1(SubCellInput2[52]), 
        .A2(SubCellInput2[53]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U2 ( .A1(SubCellInput2[55]), 
        .A2(Red_SubCellInst2_LFInst_13_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U1 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[54]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[14])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U3 ( .A1(SubCellInput2[56]), 
        .A2(SubCellInput2[57]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U2 ( .A1(SubCellInput2[59]), 
        .A2(Red_SubCellInst2_LFInst_14_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U1 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[58]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n7) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_0_n9), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_0_n8), .ZN(Red_ShiftRowsOutput2[15])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U3 ( .A1(SubCellInput2[60]), 
        .A2(SubCellInput2[61]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n8) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U2 ( .A1(SubCellInput2[63]), 
        .A2(Red_SubCellInst2_LFInst_15_LFInst_0_n7), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n9) );
  OR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U1 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[62]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_v0_0Inst_0_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_0[3]), .Z(Red_MCInst2_MC0_v0_0_0_) );
  XOR2_X1 Red_MCInst2_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_3[0]), .Z(Red_MCInst2_MC0_v0_2_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v0_3Inst_0_U2 ( .A(Red_MCInst2_MC0_v0_3Inst_0_n3), 
        .B(MCInst2_MC0_v0_3[3]), .ZN(Red_MCInst2_MC0_v0_3_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), .B(
        MCInst2_MC0_v0_0[3]), .ZN(Red_MCInst2_MC0_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U3 ( .A(Red_MCInst2_MC0_v1_0Inst_0_n6), 
        .B(Red_MCInst2_MC0_v1_0Inst_0_n5), .ZN(Red_MCInst2_MC0_v1_0_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC0_v1_1_0_), .B(
        MCInst2_MC0_v1_0[3]), .ZN(Red_MCInst2_MC0_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .Z(Red_MCInst2_MC0_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC0_v1_2Inst_0_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        Red_MCInst2_MC0_v1_1_0_), .Z(Red_MCInst2_MC0_v1_2_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v1_3Inst_0_U2 ( .A(Red_MCInst2_MC0_v1_3Inst_0_n3), 
        .B(Red_MCInst2_MC0_v1_1_0_), .ZN(Red_MCInst2_MC0_v1_3_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v1_3Inst_0_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(Red_MCInst2_MC0_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v2_0Inst_0_U2 ( .A(Red_MCInst2_MC0_v2_0Inst_0_n3), 
        .B(MCInst2_MC0_v2_0[3]), .ZN(Red_MCInst2_MC0_v2_0_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v2_0Inst_0_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .ZN(Red_MCInst2_MC0_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC0_v2_1Inst_0_U1 ( .A(MCInst2_MC0_v2_0[3]), .B(
        MCInst2_MC0_v2_0[0]), .Z(Red_MCInst2_MC0_v2_1_0_) );
  XOR2_X1 Red_MCInst2_MC0_v2_2Inst_0_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[3]), .Z(Red_MCInst2_MC0_v2_2_0_) );
  XOR2_X1 Red_MCInst2_MC0_v2_3Inst_0_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[0]), .Z(Red_MCInst2_MC0_v2_3_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v3_0Inst_0_U2 ( .A(Red_MCInst2_MC0_v3_0Inst_0_n3), 
        .B(Red_MCInst2_MC0_v3_1_0_), .ZN(Red_MCInst2_MC0_v3_0_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v3_0Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[2]), .ZN(Red_MCInst2_MC0_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U2 ( .A(Red_MCInst2_MC0_v3_2Inst_0_n3), 
        .B(MCInst2_MC0_v3_2[2]), .ZN(Red_MCInst2_MC0_v3_2_0_) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U1 ( .A(MCInst2_MC0_v3_0[2]), .B(
        Red_MCInst2_MC0_v3_1_0_), .ZN(Red_MCInst2_MC0_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC0_v3_3Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_2[2]), .Z(Red_MCInst2_MC0_v3_3_0_) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[15]) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_0_0_), 
        .B(Red_MCInst2_MC0_v1_0_0_), .ZN(Red_MCInst2_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_0_0_), 
        .B(Red_MCInst2_MC0_v3_0_0_), .Z(Red_MCInst2_MC0_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[11]) );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_1_0_), 
        .B(Red_MCInst2_MC0_v1_1_0_), .ZN(Red_MCInst2_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), 
        .B(Red_MCInst2_MC0_v3_1_0_), .Z(Red_MCInst2_MC0_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[7]) );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_2_0_), 
        .B(Red_MCInst2_MC0_v1_2_0_), .ZN(Red_MCInst2_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_2_0_), 
        .B(Red_MCInst2_MC0_v3_2_0_), .Z(Red_MCInst2_MC0_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[3]) );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_3_0_), 
        .B(Red_MCInst2_MC0_v1_3_0_), .ZN(Red_MCInst2_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_3_0_), 
        .B(Red_MCInst2_MC0_v3_3_0_), .Z(Red_MCInst2_MC0_r3Inst_XORInst_0_0_n8)
         );
  XOR2_X1 Red_MCInst2_MC1_v0_0Inst_0_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_0[3]), .Z(Red_MCInst2_MC1_v0_0_0_) );
  XOR2_X1 Red_MCInst2_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_3[0]), .Z(Red_MCInst2_MC1_v0_2_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v0_3Inst_0_U2 ( .A(Red_MCInst2_MC1_v0_3Inst_0_n3), 
        .B(MCInst2_MC1_v0_3[3]), .ZN(Red_MCInst2_MC1_v0_3_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), .B(
        MCInst2_MC1_v0_0[3]), .ZN(Red_MCInst2_MC1_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U3 ( .A(Red_MCInst2_MC1_v1_0Inst_0_n6), 
        .B(Red_MCInst2_MC1_v1_0Inst_0_n5), .ZN(Red_MCInst2_MC1_v1_0_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC1_v1_1_0_), .B(
        MCInst2_MC1_v1_0[3]), .ZN(Red_MCInst2_MC1_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .Z(Red_MCInst2_MC1_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC1_v1_2Inst_0_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        Red_MCInst2_MC1_v1_1_0_), .Z(Red_MCInst2_MC1_v1_2_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v1_3Inst_0_U2 ( .A(Red_MCInst2_MC1_v1_3Inst_0_n3), 
        .B(Red_MCInst2_MC1_v1_1_0_), .ZN(Red_MCInst2_MC1_v1_3_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v1_3Inst_0_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(Red_MCInst2_MC1_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v2_0Inst_0_U2 ( .A(Red_MCInst2_MC1_v2_0Inst_0_n3), 
        .B(MCInst2_MC1_v2_0[3]), .ZN(Red_MCInst2_MC1_v2_0_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v2_0Inst_0_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .ZN(Red_MCInst2_MC1_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC1_v2_1Inst_0_U1 ( .A(MCInst2_MC1_v2_0[3]), .B(
        MCInst2_MC1_v2_0[0]), .Z(Red_MCInst2_MC1_v2_1_0_) );
  XOR2_X1 Red_MCInst2_MC1_v2_2Inst_0_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[3]), .Z(Red_MCInst2_MC1_v2_2_0_) );
  XOR2_X1 Red_MCInst2_MC1_v2_3Inst_0_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[0]), .Z(Red_MCInst2_MC1_v2_3_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v3_0Inst_0_U2 ( .A(Red_MCInst2_MC1_v3_0Inst_0_n3), 
        .B(Red_MCInst2_MC1_v3_1_0_), .ZN(Red_MCInst2_MC1_v3_0_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v3_0Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[2]), .ZN(Red_MCInst2_MC1_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U2 ( .A(Red_MCInst2_MC1_v3_2Inst_0_n3), 
        .B(MCInst2_MC1_v3_2[2]), .ZN(Red_MCInst2_MC1_v3_2_0_) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U1 ( .A(MCInst2_MC1_v3_0[2]), .B(
        Red_MCInst2_MC1_v3_1_0_), .ZN(Red_MCInst2_MC1_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC1_v3_3Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_2[2]), .Z(Red_MCInst2_MC1_v3_3_0_) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[14]) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_0_0_), 
        .B(Red_MCInst2_MC1_v1_0_0_), .ZN(Red_MCInst2_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_0_0_), 
        .B(Red_MCInst2_MC1_v3_0_0_), .Z(Red_MCInst2_MC1_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[10]) );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_1_0_), 
        .B(Red_MCInst2_MC1_v1_1_0_), .ZN(Red_MCInst2_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), 
        .B(Red_MCInst2_MC1_v3_1_0_), .Z(Red_MCInst2_MC1_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[6]) );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_2_0_), 
        .B(Red_MCInst2_MC1_v1_2_0_), .ZN(Red_MCInst2_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_2_0_), 
        .B(Red_MCInst2_MC1_v3_2_0_), .Z(Red_MCInst2_MC1_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[2]) );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_3_0_), 
        .B(Red_MCInst2_MC1_v1_3_0_), .ZN(Red_MCInst2_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_3_0_), 
        .B(Red_MCInst2_MC1_v3_3_0_), .Z(Red_MCInst2_MC1_r3Inst_XORInst_0_0_n8)
         );
  XOR2_X1 Red_MCInst2_MC2_v0_0Inst_0_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_0[3]), .Z(Red_MCInst2_MC2_v0_0_0_) );
  XOR2_X1 Red_MCInst2_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_3[0]), .Z(Red_MCInst2_MC2_v0_2_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v0_3Inst_0_U2 ( .A(Red_MCInst2_MC2_v0_3Inst_0_n3), 
        .B(MCInst2_MC2_v0_3[3]), .ZN(Red_MCInst2_MC2_v0_3_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), .B(
        MCInst2_MC2_v0_0[3]), .ZN(Red_MCInst2_MC2_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U3 ( .A(Red_MCInst2_MC2_v1_0Inst_0_n6), 
        .B(Red_MCInst2_MC2_v1_0Inst_0_n5), .ZN(Red_MCInst2_MC2_v1_0_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC2_v1_1_0_), .B(
        MCInst2_MC2_v1_0[3]), .ZN(Red_MCInst2_MC2_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .Z(Red_MCInst2_MC2_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC2_v1_2Inst_0_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        Red_MCInst2_MC2_v1_1_0_), .Z(Red_MCInst2_MC2_v1_2_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v1_3Inst_0_U2 ( .A(Red_MCInst2_MC2_v1_3Inst_0_n3), 
        .B(Red_MCInst2_MC2_v1_1_0_), .ZN(Red_MCInst2_MC2_v1_3_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v1_3Inst_0_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(Red_MCInst2_MC2_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v2_0Inst_0_U2 ( .A(Red_MCInst2_MC2_v2_0Inst_0_n3), 
        .B(MCInst2_MC2_v2_0[3]), .ZN(Red_MCInst2_MC2_v2_0_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v2_0Inst_0_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .ZN(Red_MCInst2_MC2_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC2_v2_1Inst_0_U1 ( .A(MCInst2_MC2_v2_0[3]), .B(
        MCInst2_MC2_v2_0[0]), .Z(Red_MCInst2_MC2_v2_1_0_) );
  XOR2_X1 Red_MCInst2_MC2_v2_2Inst_0_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[3]), .Z(Red_MCInst2_MC2_v2_2_0_) );
  XOR2_X1 Red_MCInst2_MC2_v2_3Inst_0_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[0]), .Z(Red_MCInst2_MC2_v2_3_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v3_0Inst_0_U2 ( .A(Red_MCInst2_MC2_v3_0Inst_0_n3), 
        .B(Red_MCInst2_MC2_v3_1_0_), .ZN(Red_MCInst2_MC2_v3_0_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v3_0Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[2]), .ZN(Red_MCInst2_MC2_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U2 ( .A(Red_MCInst2_MC2_v3_2Inst_0_n3), 
        .B(MCInst2_MC2_v3_2[2]), .ZN(Red_MCInst2_MC2_v3_2_0_) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U1 ( .A(MCInst2_MC2_v3_0[2]), .B(
        Red_MCInst2_MC2_v3_1_0_), .ZN(Red_MCInst2_MC2_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC2_v3_3Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_2[2]), .Z(Red_MCInst2_MC2_v3_3_0_) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[13]) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_0_0_), 
        .B(Red_MCInst2_MC2_v1_0_0_), .ZN(Red_MCInst2_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_0_0_), 
        .B(Red_MCInst2_MC2_v3_0_0_), .Z(Red_MCInst2_MC2_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[9]) );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_1_0_), 
        .B(Red_MCInst2_MC2_v1_1_0_), .ZN(Red_MCInst2_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), 
        .B(Red_MCInst2_MC2_v3_1_0_), .Z(Red_MCInst2_MC2_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[5]) );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_2_0_), 
        .B(Red_MCInst2_MC2_v1_2_0_), .ZN(Red_MCInst2_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_2_0_), 
        .B(Red_MCInst2_MC2_v3_2_0_), .Z(Red_MCInst2_MC2_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[1]) );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_3_0_), 
        .B(Red_MCInst2_MC2_v1_3_0_), .ZN(Red_MCInst2_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_3_0_), 
        .B(Red_MCInst2_MC2_v3_3_0_), .Z(Red_MCInst2_MC2_r3Inst_XORInst_0_0_n8)
         );
  XOR2_X1 Red_MCInst2_MC3_v0_0Inst_0_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_0[3]), .Z(Red_MCInst2_MC3_v0_0_0_) );
  XOR2_X1 Red_MCInst2_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_3[0]), .Z(Red_MCInst2_MC3_v0_2_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v0_3Inst_0_U2 ( .A(Red_MCInst2_MC3_v0_3Inst_0_n3), 
        .B(MCInst2_MC3_v0_3[3]), .ZN(Red_MCInst2_MC3_v0_3_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), .B(
        MCInst2_MC3_v0_0[3]), .ZN(Red_MCInst2_MC3_v0_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U3 ( .A(Red_MCInst2_MC3_v1_0Inst_0_n6), 
        .B(Red_MCInst2_MC3_v1_0Inst_0_n5), .ZN(Red_MCInst2_MC3_v1_0_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC3_v1_1_0_), .B(
        MCInst2_MC3_v1_0[3]), .ZN(Red_MCInst2_MC3_v1_0Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .Z(Red_MCInst2_MC3_v1_0Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC3_v1_2Inst_0_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        Red_MCInst2_MC3_v1_1_0_), .Z(Red_MCInst2_MC3_v1_2_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v1_3Inst_0_U2 ( .A(Red_MCInst2_MC3_v1_3Inst_0_n3), 
        .B(Red_MCInst2_MC3_v1_1_0_), .ZN(Red_MCInst2_MC3_v1_3_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v1_3Inst_0_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(Red_MCInst2_MC3_v1_3Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v2_0Inst_0_U2 ( .A(Red_MCInst2_MC3_v2_0Inst_0_n3), 
        .B(MCInst2_MC3_v2_0[3]), .ZN(Red_MCInst2_MC3_v2_0_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v2_0Inst_0_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .ZN(Red_MCInst2_MC3_v2_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC3_v2_1Inst_0_U1 ( .A(MCInst2_MC3_v2_0[3]), .B(
        MCInst2_MC3_v2_0[0]), .Z(Red_MCInst2_MC3_v2_1_0_) );
  XOR2_X1 Red_MCInst2_MC3_v2_2Inst_0_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[3]), .Z(Red_MCInst2_MC3_v2_2_0_) );
  XOR2_X1 Red_MCInst2_MC3_v2_3Inst_0_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[0]), .Z(Red_MCInst2_MC3_v2_3_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v3_0Inst_0_U2 ( .A(Red_MCInst2_MC3_v3_0Inst_0_n3), 
        .B(Red_MCInst2_MC3_v3_1_0_), .ZN(Red_MCInst2_MC3_v3_0_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v3_0Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[2]), .ZN(Red_MCInst2_MC3_v3_0Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U2 ( .A(Red_MCInst2_MC3_v3_2Inst_0_n3), 
        .B(MCInst2_MC3_v3_2[2]), .ZN(Red_MCInst2_MC3_v3_2_0_) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U1 ( .A(MCInst2_MC3_v3_0[2]), .B(
        Red_MCInst2_MC3_v3_1_0_), .ZN(Red_MCInst2_MC3_v3_2Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC3_v3_3Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_2[2]), .Z(Red_MCInst2_MC3_v3_3_0_) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[12]) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_0_0_), 
        .B(Red_MCInst2_MC3_v1_0_0_), .ZN(Red_MCInst2_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_0_0_), 
        .B(Red_MCInst2_MC3_v3_0_0_), .Z(Red_MCInst2_MC3_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[8]) );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_1_0_), 
        .B(Red_MCInst2_MC3_v1_1_0_), .ZN(Red_MCInst2_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), 
        .B(Red_MCInst2_MC3_v3_1_0_), .Z(Red_MCInst2_MC3_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[4]) );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_2_0_), 
        .B(Red_MCInst2_MC3_v1_2_0_), .ZN(Red_MCInst2_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_2_0_), 
        .B(Red_MCInst2_MC3_v3_2_0_), .Z(Red_MCInst2_MC3_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[0]) );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_3_0_), 
        .B(Red_MCInst2_MC3_v1_3_0_), .ZN(Red_MCInst2_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_3_0_), 
        .B(Red_MCInst2_MC3_v3_3_0_), .Z(Red_MCInst2_MC3_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_0_LFInst_0_n6), .B(Red_KeyInst_LFInst_0_LFInst_0_n5), .ZN(Red_RoundKey[0]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U2 ( .A(Key[2]), .B(Key[3]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .Z(
        Red_KeyInst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_1_LFInst_0_n6), .B(Red_KeyInst_LFInst_1_LFInst_0_n5), .ZN(Red_RoundKey[1]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U2 ( .A(Key[6]), .B(Key[7]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .Z(
        Red_KeyInst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_2_LFInst_0_n6), .B(Red_KeyInst_LFInst_2_LFInst_0_n5), .ZN(Red_RoundKey[2]) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U2 ( .A(Key[10]), .B(Key[11]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .Z(
        Red_KeyInst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_3_LFInst_0_n6), .B(Red_KeyInst_LFInst_3_LFInst_0_n5), .ZN(Red_RoundKey[3]) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U2 ( .A(Key[14]), .B(Key[15]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .Z(
        Red_KeyInst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_4_LFInst_0_n6), .B(Red_KeyInst_LFInst_4_LFInst_0_n5), .ZN(Red_RoundKey[4]) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U2 ( .A(Key[18]), .B(Key[19]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .Z(
        Red_KeyInst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_5_LFInst_0_n6), .B(Red_KeyInst_LFInst_5_LFInst_0_n5), .ZN(Red_RoundKey[5]) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U2 ( .A(Key[22]), .B(Key[23]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .Z(
        Red_KeyInst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_6_LFInst_0_n6), .B(Red_KeyInst_LFInst_6_LFInst_0_n5), .ZN(Red_RoundKey[6]) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U2 ( .A(Key[26]), .B(Key[27]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .Z(
        Red_KeyInst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_7_LFInst_0_n6), .B(Red_KeyInst_LFInst_7_LFInst_0_n5), .ZN(Red_RoundKey[7]) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U2 ( .A(Key[30]), .B(Key[31]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .Z(
        Red_KeyInst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_8_LFInst_0_n6), .B(Red_KeyInst_LFInst_8_LFInst_0_n5), .ZN(Red_RoundKey[8]) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U2 ( .A(Key[34]), .B(Key[35]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .Z(
        Red_KeyInst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_9_LFInst_0_n6), .B(Red_KeyInst_LFInst_9_LFInst_0_n5), .ZN(Red_RoundKey[9]) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U2 ( .A(Key[38]), .B(Key[39]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .Z(
        Red_KeyInst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_10_LFInst_0_n6), .B(
        Red_KeyInst_LFInst_10_LFInst_0_n5), .ZN(Red_RoundKey[10]) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U2 ( .A(Key[42]), .B(Key[43]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .Z(
        Red_KeyInst_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_11_LFInst_0_n6), .B(
        Red_KeyInst_LFInst_11_LFInst_0_n5), .ZN(Red_RoundKey[11]) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U2 ( .A(Key[46]), .B(Key[47]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .Z(
        Red_KeyInst_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_12_LFInst_0_n6), .B(
        Red_KeyInst_LFInst_12_LFInst_0_n5), .ZN(Red_RoundKey[12]) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U2 ( .A(Key[50]), .B(Key[51]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .Z(
        Red_KeyInst_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_13_LFInst_0_n6), .B(
        Red_KeyInst_LFInst_13_LFInst_0_n5), .ZN(Red_RoundKey[13]) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U2 ( .A(Key[54]), .B(Key[55]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .Z(
        Red_KeyInst_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_14_LFInst_0_n6), .B(
        Red_KeyInst_LFInst_14_LFInst_0_n5), .ZN(Red_RoundKey[14]) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U2 ( .A(Key[58]), .B(Key[59]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .Z(
        Red_KeyInst_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U3 ( .A(
        Red_KeyInst_LFInst_15_LFInst_0_n6), .B(
        Red_KeyInst_LFInst_15_LFInst_0_n5), .ZN(Red_RoundKey[15]) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U2 ( .A(Key[62]), .B(Key[63]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_0_n5) );
  XOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .Z(
        Red_KeyInst_LFInst_15_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_0_LFInst_0_n5), .ZN(Red_SignaltoCheck[0]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U2 ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[3]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[1]), .Z(Red_ToCheckInst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_1_LFInst_0_n5), .ZN(Red_SignaltoCheck[1]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U2 ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[7]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[5]), .Z(Red_ToCheckInst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_2_LFInst_0_n5), .ZN(Red_SignaltoCheck[2]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U2 ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[11]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[9]), .Z(Red_ToCheckInst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_3_LFInst_0_n5), .ZN(Red_SignaltoCheck[3]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U2 ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[15]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .Z(Red_ToCheckInst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_4_LFInst_0_n5), .ZN(Red_SignaltoCheck[4]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U2 ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[19]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .Z(Red_ToCheckInst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_5_LFInst_0_n5), .ZN(Red_SignaltoCheck[5]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U2 ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[23]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .Z(Red_ToCheckInst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_6_LFInst_0_n5), .ZN(Red_SignaltoCheck[6]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U2 ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[27]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .Z(Red_ToCheckInst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_7_LFInst_0_n5), .ZN(Red_SignaltoCheck[7]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U2 ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[31]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .Z(Red_ToCheckInst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_8_LFInst_0_n5), .ZN(Red_SignaltoCheck[8]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U2 ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[35]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .Z(Red_ToCheckInst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_9_LFInst_0_n5), .ZN(Red_SignaltoCheck[9]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U2 ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[39]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .Z(Red_ToCheckInst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_10_LFInst_0_n5), .ZN(Red_SignaltoCheck[10]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U2 ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[43]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .Z(Red_ToCheckInst_LFInst_10_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_11_LFInst_0_n5), .ZN(Red_SignaltoCheck[11]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U2 ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[47]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .Z(Red_ToCheckInst_LFInst_11_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_12_LFInst_0_n5), .ZN(Red_SignaltoCheck[12]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U2 ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[51]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .Z(Red_ToCheckInst_LFInst_12_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_13_LFInst_0_n5), .ZN(Red_SignaltoCheck[13]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U2 ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[55]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .Z(Red_ToCheckInst_LFInst_13_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_14_LFInst_0_n5), .ZN(Red_SignaltoCheck[14]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U2 ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[59]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .Z(Red_ToCheckInst_LFInst_14_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_15_LFInst_0_n5), .ZN(Red_SignaltoCheck[15]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U2 ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[63]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .Z(Red_ToCheckInst_LFInst_15_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_16_LFInst_0_n5), .ZN(Red_SignaltoCheck[16]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U2 ( .A(Ciphertext[2]), .B(
        Ciphertext[3]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U1 ( .A(Ciphertext[0]), .B(
        Ciphertext[1]), .Z(Red_ToCheckInst_LFInst_16_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_17_LFInst_0_n5), .ZN(Red_SignaltoCheck[17]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U2 ( .A(Ciphertext[6]), .B(
        Ciphertext[7]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U1 ( .A(Ciphertext[4]), .B(
        Ciphertext[5]), .Z(Red_ToCheckInst_LFInst_17_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_18_LFInst_0_n5), .ZN(Red_SignaltoCheck[18]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U2 ( .A(Ciphertext[10]), .B(
        Ciphertext[11]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U1 ( .A(Ciphertext[8]), .B(
        Ciphertext[9]), .Z(Red_ToCheckInst_LFInst_18_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_19_LFInst_0_n5), .ZN(Red_SignaltoCheck[19]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U2 ( .A(Ciphertext[14]), .B(
        Ciphertext[15]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U1 ( .A(Ciphertext[12]), .B(
        Ciphertext[13]), .Z(Red_ToCheckInst_LFInst_19_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_20_LFInst_0_n5), .ZN(Red_SignaltoCheck[20]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U2 ( .A(Ciphertext[18]), .B(
        Ciphertext[19]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U1 ( .A(Ciphertext[16]), .B(
        Ciphertext[17]), .Z(Red_ToCheckInst_LFInst_20_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_21_LFInst_0_n5), .ZN(Red_SignaltoCheck[21]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U2 ( .A(Ciphertext[22]), .B(
        Ciphertext[23]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U1 ( .A(Ciphertext[20]), .B(
        Ciphertext[21]), .Z(Red_ToCheckInst_LFInst_21_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_22_LFInst_0_n5), .ZN(Red_SignaltoCheck[22]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U2 ( .A(Ciphertext[26]), .B(
        Ciphertext[27]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U1 ( .A(Ciphertext[24]), .B(
        Ciphertext[25]), .Z(Red_ToCheckInst_LFInst_22_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_23_LFInst_0_n5), .ZN(Red_SignaltoCheck[23]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U2 ( .A(Ciphertext[30]), .B(
        Ciphertext[31]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U1 ( .A(Ciphertext[28]), .B(
        Ciphertext[29]), .Z(Red_ToCheckInst_LFInst_23_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_24_LFInst_0_n5), .ZN(Red_SignaltoCheck[24]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U2 ( .A(Ciphertext[34]), .B(
        Ciphertext[35]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U1 ( .A(Ciphertext[32]), .B(
        Ciphertext[33]), .Z(Red_ToCheckInst_LFInst_24_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_25_LFInst_0_n5), .ZN(Red_SignaltoCheck[25]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U2 ( .A(Ciphertext[38]), .B(
        Ciphertext[39]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U1 ( .A(Ciphertext[36]), .B(
        Ciphertext[37]), .Z(Red_ToCheckInst_LFInst_25_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_26_LFInst_0_n5), .ZN(Red_SignaltoCheck[26]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U2 ( .A(Ciphertext[42]), .B(
        Ciphertext[43]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U1 ( .A(Ciphertext[40]), .B(
        Ciphertext[41]), .Z(Red_ToCheckInst_LFInst_26_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_27_LFInst_0_n5), .ZN(Red_SignaltoCheck[27]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U2 ( .A(Ciphertext[46]), .B(
        Ciphertext[47]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U1 ( .A(Ciphertext[44]), .B(
        Ciphertext[45]), .Z(Red_ToCheckInst_LFInst_27_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_28_LFInst_0_n5), .ZN(Red_SignaltoCheck[28]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U2 ( .A(Ciphertext[50]), .B(
        Ciphertext[51]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U1 ( .A(Ciphertext[48]), .B(
        Ciphertext[49]), .Z(Red_ToCheckInst_LFInst_28_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_29_LFInst_0_n5), .ZN(Red_SignaltoCheck[29]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U2 ( .A(Ciphertext[54]), .B(
        Ciphertext[55]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U1 ( .A(Ciphertext[52]), .B(
        Ciphertext[53]), .Z(Red_ToCheckInst_LFInst_29_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_30_LFInst_0_n5), .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U2 ( .A(Ciphertext[58]), .B(
        Ciphertext[59]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U1 ( .A(Ciphertext[56]), .B(
        Ciphertext[57]), .Z(Red_ToCheckInst_LFInst_30_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_31_LFInst_0_n5), .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U2 ( .A(Ciphertext[62]), .B(
        Ciphertext[63]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U1 ( .A(Ciphertext[60]), .B(
        Ciphertext[61]), .Z(Red_ToCheckInst_LFInst_31_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_32_LFInst_0_n5), .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U2 ( .A(Red_MCInst2_MC3_v3_1_0_), 
        .B(MCInst2_MC3_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[2]), .Z(Red_ToCheckInst_LFInst_32_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_33_LFInst_0_n5), .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U2 ( .A(Red_MCInst2_MC2_v3_1_0_), 
        .B(MCInst2_MC2_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[2]), .Z(Red_ToCheckInst_LFInst_33_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_34_LFInst_0_n5), .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U2 ( .A(Red_MCInst2_MC1_v3_1_0_), 
        .B(MCInst2_MC1_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[2]), .Z(Red_ToCheckInst_LFInst_34_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_35_LFInst_0_n5), .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U2 ( .A(Red_MCInst2_MC0_v3_1_0_), 
        .B(MCInst2_MC0_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[2]), .Z(Red_ToCheckInst_LFInst_35_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_36_LFInst_0_n5), .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U2 ( .A(MCInst2_MC3_v2_0[3]), 
        .B(MCInst2_MC3_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(Red_ToCheckInst_LFInst_36_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_37_LFInst_0_n5), .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U2 ( .A(MCInst2_MC2_v2_0[3]), 
        .B(MCInst2_MC2_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(Red_ToCheckInst_LFInst_37_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_38_LFInst_0_n5), .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U2 ( .A(MCInst2_MC1_v2_0[3]), 
        .B(MCInst2_MC1_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(Red_ToCheckInst_LFInst_38_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_39_LFInst_0_n5), .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U2 ( .A(MCInst2_MC0_v2_0[3]), 
        .B(MCInst2_MC0_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(Red_ToCheckInst_LFInst_39_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_40_LFInst_0_n5), .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U2 ( .A(Red_MCInst2_MC3_v1_1_0_), 
        .B(MCInst2_MC3_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U1 ( .A(MCInst2_MC3_v1_0[0]), .B(
        MCInst2_MC3_v1_3[2]), .Z(Red_ToCheckInst_LFInst_40_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_41_LFInst_0_n5), .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U2 ( .A(Red_MCInst2_MC2_v1_1_0_), 
        .B(MCInst2_MC2_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U1 ( .A(MCInst2_MC2_v1_0[0]), .B(
        MCInst2_MC2_v1_3[2]), .Z(Red_ToCheckInst_LFInst_41_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_42_LFInst_0_n5), .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U2 ( .A(Red_MCInst2_MC1_v1_1_0_), 
        .B(MCInst2_MC1_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U1 ( .A(MCInst2_MC1_v1_0[0]), .B(
        MCInst2_MC1_v1_3[2]), .Z(Red_ToCheckInst_LFInst_42_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_43_LFInst_0_n5), .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U2 ( .A(Red_MCInst2_MC0_v1_1_0_), 
        .B(MCInst2_MC0_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U1 ( .A(MCInst2_MC0_v1_0[0]), .B(
        MCInst2_MC0_v1_3[2]), .Z(Red_ToCheckInst_LFInst_43_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_44_LFInst_0_n5), .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U2 ( .A(MCInst2_MC3_v0_3[3]), 
        .B(MCInst2_MC3_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U1 ( .A(Red_MCInst2_MC3_v0_1_0_), 
        .B(MCInst2_MC3_v0_0[3]), .Z(Red_ToCheckInst_LFInst_44_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_45_LFInst_0_n5), .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U2 ( .A(MCInst2_MC2_v0_3[3]), 
        .B(MCInst2_MC2_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U1 ( .A(Red_MCInst2_MC2_v0_1_0_), 
        .B(MCInst2_MC2_v0_0[3]), .Z(Red_ToCheckInst_LFInst_45_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_46_LFInst_0_n5), .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U2 ( .A(MCInst2_MC1_v0_3[3]), 
        .B(MCInst2_MC1_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U1 ( .A(Red_MCInst2_MC1_v0_1_0_), 
        .B(MCInst2_MC1_v0_0[3]), .Z(Red_ToCheckInst_LFInst_46_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_47_LFInst_0_n5), .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U2 ( .A(MCInst2_MC0_v0_3[3]), 
        .B(MCInst2_MC0_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U1 ( .A(Red_MCInst2_MC0_v0_1_0_), 
        .B(MCInst2_MC0_v0_0[3]), .Z(Red_ToCheckInst_LFInst_47_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_48_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_48_LFInst_0_n5), .ZN(Red_SignaltoCheck[48]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U2 ( .A(SubCellInput2[2]), .B(
        SubCellInput2[3]), .ZN(Red_ToCheckInst_LFInst_48_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U1 ( .A(SubCellInput2[0]), .B(
        SubCellInput2[1]), .Z(Red_ToCheckInst_LFInst_48_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_49_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_49_LFInst_0_n5), .ZN(Red_SignaltoCheck[49]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U2 ( .A(SubCellInput2[6]), .B(
        SubCellInput2[7]), .ZN(Red_ToCheckInst_LFInst_49_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U1 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[5]), .Z(Red_ToCheckInst_LFInst_49_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_50_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_50_LFInst_0_n5), .ZN(Red_SignaltoCheck[50]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U2 ( .A(SubCellInput2[10]), .B(
        SubCellInput2[11]), .ZN(Red_ToCheckInst_LFInst_50_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U1 ( .A(SubCellInput2[8]), .B(
        SubCellInput2[9]), .Z(Red_ToCheckInst_LFInst_50_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_51_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_51_LFInst_0_n5), .ZN(Red_SignaltoCheck[51]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U2 ( .A(SubCellInput2[14]), .B(
        SubCellInput2[15]), .ZN(Red_ToCheckInst_LFInst_51_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U1 ( .A(SubCellInput2[12]), .B(
        SubCellInput2[13]), .Z(Red_ToCheckInst_LFInst_51_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_52_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_52_LFInst_0_n5), .ZN(Red_SignaltoCheck[52]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U2 ( .A(SubCellInput2[18]), .B(
        SubCellInput2[19]), .ZN(Red_ToCheckInst_LFInst_52_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U1 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[17]), .Z(Red_ToCheckInst_LFInst_52_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_53_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_53_LFInst_0_n5), .ZN(Red_SignaltoCheck[53]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U2 ( .A(SubCellInput2[22]), .B(
        SubCellInput2[23]), .ZN(Red_ToCheckInst_LFInst_53_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U1 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[21]), .Z(Red_ToCheckInst_LFInst_53_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_54_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_54_LFInst_0_n5), .ZN(Red_SignaltoCheck[54]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U2 ( .A(SubCellInput2[26]), .B(
        SubCellInput2[27]), .ZN(Red_ToCheckInst_LFInst_54_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U1 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[25]), .Z(Red_ToCheckInst_LFInst_54_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_55_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_55_LFInst_0_n5), .ZN(Red_SignaltoCheck[55]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U2 ( .A(SubCellInput2[30]), .B(
        SubCellInput2[31]), .ZN(Red_ToCheckInst_LFInst_55_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U1 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[29]), .Z(Red_ToCheckInst_LFInst_55_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_56_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_56_LFInst_0_n5), .ZN(Red_SignaltoCheck[56]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U2 ( .A(SubCellInput2[34]), .B(
        SubCellInput2[35]), .ZN(Red_ToCheckInst_LFInst_56_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U1 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[33]), .Z(Red_ToCheckInst_LFInst_56_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_57_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_57_LFInst_0_n5), .ZN(Red_SignaltoCheck[57]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U2 ( .A(SubCellInput2[38]), .B(
        SubCellInput2[39]), .ZN(Red_ToCheckInst_LFInst_57_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U1 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[37]), .Z(Red_ToCheckInst_LFInst_57_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_58_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_58_LFInst_0_n5), .ZN(Red_SignaltoCheck[58]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U2 ( .A(SubCellInput2[42]), .B(
        SubCellInput2[43]), .ZN(Red_ToCheckInst_LFInst_58_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U1 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[41]), .Z(Red_ToCheckInst_LFInst_58_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_59_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_59_LFInst_0_n5), .ZN(Red_SignaltoCheck[59]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U2 ( .A(SubCellInput2[46]), .B(
        SubCellInput2[47]), .ZN(Red_ToCheckInst_LFInst_59_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U1 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[45]), .Z(Red_ToCheckInst_LFInst_59_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_60_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_60_LFInst_0_n5), .ZN(Red_SignaltoCheck[60]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U2 ( .A(SubCellInput2[50]), .B(
        SubCellInput2[51]), .ZN(Red_ToCheckInst_LFInst_60_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U1 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[49]), .Z(Red_ToCheckInst_LFInst_60_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_61_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_61_LFInst_0_n5), .ZN(Red_SignaltoCheck[61]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U2 ( .A(SubCellInput2[54]), .B(
        SubCellInput2[55]), .ZN(Red_ToCheckInst_LFInst_61_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U1 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[53]), .Z(Red_ToCheckInst_LFInst_61_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_62_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_62_LFInst_0_n5), .ZN(Red_SignaltoCheck[62]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U2 ( .A(SubCellInput2[58]), .B(
        SubCellInput2[59]), .ZN(Red_ToCheckInst_LFInst_62_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U1 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[57]), .Z(Red_ToCheckInst_LFInst_62_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_63_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_63_LFInst_0_n5), .ZN(Red_SignaltoCheck[63]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U2 ( .A(SubCellInput2[62]), .B(
        SubCellInput2[63]), .ZN(Red_ToCheckInst_LFInst_63_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U1 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[61]), .Z(Red_ToCheckInst_LFInst_63_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_64_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_64_LFInst_0_n5), .ZN(Red_SignaltoCheck[64]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U2 ( .A(MC_output[2]), .B(
        MC_output[3]), .ZN(Red_ToCheckInst_LFInst_64_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U1 ( .A(MC_output[0]), .B(
        MC_output[1]), .Z(Red_ToCheckInst_LFInst_64_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_65_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_65_LFInst_0_n5), .ZN(Red_SignaltoCheck[65]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U2 ( .A(MC_output[6]), .B(
        MC_output[7]), .ZN(Red_ToCheckInst_LFInst_65_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U1 ( .A(MC_output[4]), .B(
        MC_output[5]), .Z(Red_ToCheckInst_LFInst_65_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_66_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_66_LFInst_0_n5), .ZN(Red_SignaltoCheck[66]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U2 ( .A(MC_output[10]), .B(
        MC_output[11]), .ZN(Red_ToCheckInst_LFInst_66_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U1 ( .A(MC_output[8]), .B(
        MC_output[9]), .Z(Red_ToCheckInst_LFInst_66_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_67_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_67_LFInst_0_n5), .ZN(Red_SignaltoCheck[67]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U2 ( .A(MC_output[14]), .B(
        MC_output[15]), .ZN(Red_ToCheckInst_LFInst_67_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U1 ( .A(MC_output[12]), .B(
        MC_output[13]), .Z(Red_ToCheckInst_LFInst_67_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_68_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_68_LFInst_0_n5), .ZN(Red_SignaltoCheck[68]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U2 ( .A(MC_output[18]), .B(
        MC_output[19]), .ZN(Red_ToCheckInst_LFInst_68_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U1 ( .A(MC_output[16]), .B(
        MC_output[17]), .Z(Red_ToCheckInst_LFInst_68_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_69_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_69_LFInst_0_n5), .ZN(Red_SignaltoCheck[69]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U2 ( .A(MC_output[22]), .B(
        MC_output[23]), .ZN(Red_ToCheckInst_LFInst_69_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U1 ( .A(MC_output[20]), .B(
        MC_output[21]), .Z(Red_ToCheckInst_LFInst_69_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_70_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_70_LFInst_0_n5), .ZN(Red_SignaltoCheck[70]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U2 ( .A(MC_output[26]), .B(
        MC_output[27]), .ZN(Red_ToCheckInst_LFInst_70_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U1 ( .A(MC_output[24]), .B(
        MC_output[25]), .Z(Red_ToCheckInst_LFInst_70_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_71_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_71_LFInst_0_n5), .ZN(Red_SignaltoCheck[71]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U2 ( .A(MC_output[30]), .B(
        MC_output[31]), .ZN(Red_ToCheckInst_LFInst_71_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U1 ( .A(MC_output[28]), .B(
        MC_output[29]), .Z(Red_ToCheckInst_LFInst_71_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_72_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_72_LFInst_0_n5), .ZN(Red_SignaltoCheck[72]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U2 ( .A(MC_output[34]), .B(
        MC_output[35]), .ZN(Red_ToCheckInst_LFInst_72_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U1 ( .A(MC_output[32]), .B(
        MC_output[33]), .Z(Red_ToCheckInst_LFInst_72_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_73_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_73_LFInst_0_n5), .ZN(Red_SignaltoCheck[73]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U2 ( .A(MC_output[38]), .B(
        MC_output[39]), .ZN(Red_ToCheckInst_LFInst_73_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U1 ( .A(MC_output[36]), .B(
        MC_output[37]), .Z(Red_ToCheckInst_LFInst_73_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_74_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_74_LFInst_0_n5), .ZN(Red_SignaltoCheck[74]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U2 ( .A(MC_output[42]), .B(
        MC_output[43]), .ZN(Red_ToCheckInst_LFInst_74_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U1 ( .A(MC_output[40]), .B(
        MC_output[41]), .Z(Red_ToCheckInst_LFInst_74_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_75_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_75_LFInst_0_n5), .ZN(Red_SignaltoCheck[75]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U2 ( .A(MC_output[46]), .B(
        MC_output[47]), .ZN(Red_ToCheckInst_LFInst_75_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U1 ( .A(MC_output[44]), .B(
        MC_output[45]), .Z(Red_ToCheckInst_LFInst_75_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_76_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_76_LFInst_0_n5), .ZN(Red_SignaltoCheck[76]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U2 ( .A(MC_output[50]), .B(
        MC_output[51]), .ZN(Red_ToCheckInst_LFInst_76_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U1 ( .A(MC_output[48]), .B(
        MC_output[49]), .Z(Red_ToCheckInst_LFInst_76_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_77_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_77_LFInst_0_n5), .ZN(Red_SignaltoCheck[77]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U2 ( .A(MC_output[54]), .B(
        MC_output[55]), .ZN(Red_ToCheckInst_LFInst_77_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U1 ( .A(MC_output[52]), .B(
        MC_output[53]), .Z(Red_ToCheckInst_LFInst_77_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_78_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_78_LFInst_0_n5), .ZN(Red_SignaltoCheck[78]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U2 ( .A(MC_output[58]), .B(
        MC_output[59]), .ZN(Red_ToCheckInst_LFInst_78_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U1 ( .A(MC_output[56]), .B(
        MC_output[57]), .Z(Red_ToCheckInst_LFInst_78_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_79_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_79_LFInst_0_n5), .ZN(Red_SignaltoCheck[79]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U2 ( .A(MC_output[62]), .B(
        MC_output[63]), .ZN(Red_ToCheckInst_LFInst_79_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U1 ( .A(MC_output[60]), .B(
        MC_output[61]), .Z(Red_ToCheckInst_LFInst_79_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_80_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_80_LFInst_0_n5), .ZN(Red_SignaltoCheck[80]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U2 ( .A(Red_MCInst_MC3_v3_1_0_), 
        .B(MCInst_MC3_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_80_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[2]), .Z(Red_ToCheckInst_LFInst_80_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_81_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_81_LFInst_0_n5), .ZN(Red_SignaltoCheck[81]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U2 ( .A(Red_MCInst_MC2_v3_1_0_), 
        .B(MCInst_MC2_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_81_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[2]), .Z(Red_ToCheckInst_LFInst_81_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_82_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_82_LFInst_0_n5), .ZN(Red_SignaltoCheck[82]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U2 ( .A(Red_MCInst_MC1_v3_1_0_), 
        .B(MCInst_MC1_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_82_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[2]), .Z(Red_ToCheckInst_LFInst_82_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_83_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_83_LFInst_0_n5), .ZN(Red_SignaltoCheck[83]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U2 ( .A(Red_MCInst_MC0_v3_1_0_), 
        .B(MCInst_MC0_v3_2[2]), .ZN(Red_ToCheckInst_LFInst_83_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[2]), .Z(Red_ToCheckInst_LFInst_83_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_84_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_84_LFInst_0_n5), .ZN(Red_SignaltoCheck[84]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        MCInst_MC3_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_84_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(Red_ToCheckInst_LFInst_84_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_85_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_85_LFInst_0_n5), .ZN(Red_SignaltoCheck[85]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        MCInst_MC2_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_85_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(Red_ToCheckInst_LFInst_85_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_86_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_86_LFInst_0_n5), .ZN(Red_SignaltoCheck[86]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        MCInst_MC1_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_86_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(Red_ToCheckInst_LFInst_86_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_87_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_87_LFInst_0_n5), .ZN(Red_SignaltoCheck[87]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        MCInst_MC0_v2_0[0]), .ZN(Red_ToCheckInst_LFInst_87_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(Red_ToCheckInst_LFInst_87_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_88_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_88_LFInst_0_n5), .ZN(Red_SignaltoCheck[88]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U2 ( .A(Red_MCInst_MC3_v1_1_0_), 
        .B(MCInst_MC3_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_88_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U1 ( .A(MCInst_MC3_v1_0[0]), .B(
        MCInst_MC3_v1_3[2]), .Z(Red_ToCheckInst_LFInst_88_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_89_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_89_LFInst_0_n5), .ZN(Red_SignaltoCheck[89]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U2 ( .A(Red_MCInst_MC2_v1_1_0_), 
        .B(MCInst_MC2_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_89_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U1 ( .A(MCInst_MC2_v1_0[0]), .B(
        MCInst_MC2_v1_3[2]), .Z(Red_ToCheckInst_LFInst_89_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_90_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_90_LFInst_0_n5), .ZN(Red_SignaltoCheck[90]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U2 ( .A(Red_MCInst_MC1_v1_1_0_), 
        .B(MCInst_MC1_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_90_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U1 ( .A(MCInst_MC1_v1_0[0]), .B(
        MCInst_MC1_v1_3[2]), .Z(Red_ToCheckInst_LFInst_90_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_91_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_91_LFInst_0_n5), .ZN(Red_SignaltoCheck[91]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U2 ( .A(Red_MCInst_MC0_v1_1_0_), 
        .B(MCInst_MC0_v1_0[3]), .ZN(Red_ToCheckInst_LFInst_91_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U1 ( .A(MCInst_MC0_v1_0[0]), .B(
        MCInst_MC0_v1_3[2]), .Z(Red_ToCheckInst_LFInst_91_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_92_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_92_LFInst_0_n5), .ZN(Red_SignaltoCheck[92]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U2 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_92_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U1 ( .A(Red_MCInst_MC3_v0_1_0_), 
        .B(MCInst_MC3_v0_0[3]), .Z(Red_ToCheckInst_LFInst_92_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_93_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_93_LFInst_0_n5), .ZN(Red_SignaltoCheck[93]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U2 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_93_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U1 ( .A(Red_MCInst_MC2_v0_1_0_), 
        .B(MCInst_MC2_v0_0[3]), .Z(Red_ToCheckInst_LFInst_93_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_94_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_94_LFInst_0_n5), .ZN(Red_SignaltoCheck[94]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U2 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_94_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U1 ( .A(Red_MCInst_MC1_v0_1_0_), 
        .B(MCInst_MC1_v0_0[3]), .Z(Red_ToCheckInst_LFInst_94_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_95_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_95_LFInst_0_n5), .ZN(Red_SignaltoCheck[95]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U2 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v0_3[0]), .ZN(Red_ToCheckInst_LFInst_95_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U1 ( .A(Red_MCInst_MC0_v0_1_0_), 
        .B(MCInst_MC0_v0_0[3]), .Z(Red_ToCheckInst_LFInst_95_LFInst_0_n6) );
  NOR2_X1 Check1_CheckInst_0_U191 ( .A1(Check1_CheckInst_0_n190), .A2(
        Check1_CheckInst_0_n189), .ZN(Error_0_) );
  NAND2_X1 Check1_CheckInst_0_U190 ( .A1(Check1_CheckInst_0_n188), .A2(
        Check1_CheckInst_0_n187), .ZN(Check1_CheckInst_0_n189) );
  NOR2_X1 Check1_CheckInst_0_U189 ( .A1(Check1_CheckInst_0_n186), .A2(
        Check1_CheckInst_0_n185), .ZN(Check1_CheckInst_0_n187) );
  NAND2_X1 Check1_CheckInst_0_U188 ( .A1(Check1_CheckInst_0_n184), .A2(
        Check1_CheckInst_0_n183), .ZN(Check1_CheckInst_0_n185) );
  NOR2_X1 Check1_CheckInst_0_U187 ( .A1(Check1_CheckInst_0_n182), .A2(
        Check1_CheckInst_0_n181), .ZN(Check1_CheckInst_0_n183) );
  NAND2_X1 Check1_CheckInst_0_U186 ( .A1(Check1_CheckInst_0_n180), .A2(
        Check1_CheckInst_0_n179), .ZN(Check1_CheckInst_0_n181) );
  NOR2_X1 Check1_CheckInst_0_U185 ( .A1(Check1_CheckInst_0_n178), .A2(
        Check1_CheckInst_0_n177), .ZN(Check1_CheckInst_0_n179) );
  NAND2_X1 Check1_CheckInst_0_U184 ( .A1(Check1_CheckInst_0_n176), .A2(
        Check1_CheckInst_0_n175), .ZN(Check1_CheckInst_0_n177) );
  NOR2_X1 Check1_CheckInst_0_U183 ( .A1(Check1_CheckInst_0_n174), .A2(
        Check1_CheckInst_0_n173), .ZN(Check1_CheckInst_0_n175) );
  NAND2_X1 Check1_CheckInst_0_U182 ( .A1(Check1_CheckInst_0_n172), .A2(
        Check1_CheckInst_0_n171), .ZN(Check1_CheckInst_0_n173) );
  XNOR2_X1 Check1_CheckInst_0_U181 ( .A(Red_ShiftRowsOutput[10]), .B(
        Red_SignaltoCheck[90]), .ZN(Check1_CheckInst_0_n171) );
  XNOR2_X1 Check1_CheckInst_0_U180 ( .A(Red_ShiftRowsOutput[12]), .B(
        Red_SignaltoCheck[92]), .ZN(Check1_CheckInst_0_n172) );
  NAND2_X1 Check1_CheckInst_0_U179 ( .A1(Check1_CheckInst_0_n170), .A2(
        Check1_CheckInst_0_n169), .ZN(Check1_CheckInst_0_n174) );
  XNOR2_X1 Check1_CheckInst_0_U178 ( .A(Red_ShiftRowsOutput[9]), .B(
        Red_SignaltoCheck[89]), .ZN(Check1_CheckInst_0_n169) );
  XNOR2_X1 Check1_CheckInst_0_U177 ( .A(Red_ShiftRowsOutput[11]), .B(
        Red_SignaltoCheck[91]), .ZN(Check1_CheckInst_0_n170) );
  NOR2_X1 Check1_CheckInst_0_U176 ( .A1(Check1_CheckInst_0_n168), .A2(
        Check1_CheckInst_0_n167), .ZN(Check1_CheckInst_0_n176) );
  XOR2_X1 Check1_CheckInst_0_U175 ( .A(Red_MC_output[12]), .B(
        Red_SignaltoCheck[76]), .Z(Check1_CheckInst_0_n167) );
  XOR2_X1 Check1_CheckInst_0_U174 ( .A(Red_MC_output[11]), .B(
        Red_SignaltoCheck[75]), .Z(Check1_CheckInst_0_n168) );
  NAND2_X1 Check1_CheckInst_0_U173 ( .A1(Check1_CheckInst_0_n166), .A2(
        Check1_CheckInst_0_n165), .ZN(Check1_CheckInst_0_n178) );
  XNOR2_X1 Check1_CheckInst_0_U172 ( .A(Red_MC_output[8]), .B(
        Red_SignaltoCheck[72]), .ZN(Check1_CheckInst_0_n165) );
  XNOR2_X1 Check1_CheckInst_0_U171 ( .A(Red_MC_output[10]), .B(
        Red_SignaltoCheck[74]), .ZN(Check1_CheckInst_0_n166) );
  NOR2_X1 Check1_CheckInst_0_U170 ( .A1(Check1_CheckInst_0_n164), .A2(
        Check1_CheckInst_0_n163), .ZN(Check1_CheckInst_0_n180) );
  NAND2_X1 Check1_CheckInst_0_U169 ( .A1(Check1_CheckInst_0_n162), .A2(
        Check1_CheckInst_0_n161), .ZN(Check1_CheckInst_0_n163) );
  NOR2_X1 Check1_CheckInst_0_U168 ( .A1(Check1_CheckInst_0_n160), .A2(
        Check1_CheckInst_0_n159), .ZN(Check1_CheckInst_0_n161) );
  NAND2_X1 Check1_CheckInst_0_U167 ( .A1(Check1_CheckInst_0_n158), .A2(
        Check1_CheckInst_0_n157), .ZN(Check1_CheckInst_0_n159) );
  XNOR2_X1 Check1_CheckInst_0_U166 ( .A(Red_MC_output[7]), .B(
        Red_SignaltoCheck[71]), .ZN(Check1_CheckInst_0_n157) );
  XNOR2_X1 Check1_CheckInst_0_U165 ( .A(Red_MC_output[9]), .B(
        Red_SignaltoCheck[73]), .ZN(Check1_CheckInst_0_n158) );
  NAND2_X1 Check1_CheckInst_0_U164 ( .A1(Check1_CheckInst_0_n156), .A2(
        Check1_CheckInst_0_n155), .ZN(Check1_CheckInst_0_n160) );
  XNOR2_X1 Check1_CheckInst_0_U163 ( .A(Red_ShiftRowsOutput[2]), .B(
        Red_SignaltoCheck[82]), .ZN(Check1_CheckInst_0_n155) );
  XNOR2_X1 Check1_CheckInst_0_U162 ( .A(Red_ShiftRowsOutput[1]), .B(
        Red_SignaltoCheck[81]), .ZN(Check1_CheckInst_0_n156) );
  NOR2_X1 Check1_CheckInst_0_U161 ( .A1(Check1_CheckInst_0_n154), .A2(
        Check1_CheckInst_0_n153), .ZN(Check1_CheckInst_0_n162) );
  XOR2_X1 Check1_CheckInst_0_U160 ( .A(Red_MC_output[14]), .B(
        Red_SignaltoCheck[78]), .Z(Check1_CheckInst_0_n153) );
  XOR2_X1 Check1_CheckInst_0_U159 ( .A(Red_ShiftRowsOutput[0]), .B(
        Red_SignaltoCheck[80]), .Z(Check1_CheckInst_0_n154) );
  NAND2_X1 Check1_CheckInst_0_U158 ( .A1(Check1_CheckInst_0_n152), .A2(
        Check1_CheckInst_0_n151), .ZN(Check1_CheckInst_0_n164) );
  XNOR2_X1 Check1_CheckInst_0_U157 ( .A(Red_MC_output[13]), .B(
        Red_SignaltoCheck[77]), .ZN(Check1_CheckInst_0_n151) );
  XNOR2_X1 Check1_CheckInst_0_U156 ( .A(Red_MC_output[15]), .B(
        Red_SignaltoCheck[79]), .ZN(Check1_CheckInst_0_n152) );
  NAND2_X1 Check1_CheckInst_0_U155 ( .A1(Check1_CheckInst_0_n150), .A2(
        Check1_CheckInst_0_n149), .ZN(Check1_CheckInst_0_n182) );
  NOR2_X1 Check1_CheckInst_0_U154 ( .A1(Check1_CheckInst_0_n148), .A2(
        Check1_CheckInst_0_n147), .ZN(Check1_CheckInst_0_n149) );
  NAND2_X1 Check1_CheckInst_0_U153 ( .A1(Check1_CheckInst_0_n146), .A2(
        Check1_CheckInst_0_n145), .ZN(Check1_CheckInst_0_n147) );
  NOR2_X1 Check1_CheckInst_0_U152 ( .A1(Check1_CheckInst_0_n144), .A2(
        Check1_CheckInst_0_n143), .ZN(Check1_CheckInst_0_n145) );
  XOR2_X1 Check1_CheckInst_0_U151 ( .A(Red_MC_output2[15]), .B(
        Red_SignaltoCheck[31]), .Z(Check1_CheckInst_0_n143) );
  XOR2_X1 Check1_CheckInst_0_U150 ( .A(Red_MC_output2[14]), .B(
        Red_SignaltoCheck[30]), .Z(Check1_CheckInst_0_n144) );
  NOR2_X1 Check1_CheckInst_0_U149 ( .A1(Check1_CheckInst_0_n142), .A2(
        Check1_CheckInst_0_n141), .ZN(Check1_CheckInst_0_n146) );
  XOR2_X1 Check1_CheckInst_0_U148 ( .A(Red_ShiftRowsOutput2[1]), .B(
        Red_SignaltoCheck[33]), .Z(Check1_CheckInst_0_n141) );
  XOR2_X1 Check1_CheckInst_0_U147 ( .A(Red_MC_output2[13]), .B(
        Red_SignaltoCheck[29]), .Z(Check1_CheckInst_0_n142) );
  NAND2_X1 Check1_CheckInst_0_U146 ( .A1(Check1_CheckInst_0_n140), .A2(
        Check1_CheckInst_0_n139), .ZN(Check1_CheckInst_0_n148) );
  XNOR2_X1 Check1_CheckInst_0_U145 ( .A(Red_ShiftRowsOutput2[0]), .B(
        Red_SignaltoCheck[32]), .ZN(Check1_CheckInst_0_n139) );
  XNOR2_X1 Check1_CheckInst_0_U144 ( .A(Red_ShiftRowsOutput2[2]), .B(
        Red_SignaltoCheck[34]), .ZN(Check1_CheckInst_0_n140) );
  NOR2_X1 Check1_CheckInst_0_U143 ( .A1(Check1_CheckInst_0_n138), .A2(
        Check1_CheckInst_0_n137), .ZN(Check1_CheckInst_0_n150) );
  XOR2_X1 Check1_CheckInst_0_U142 ( .A(Red_MC_output2[9]), .B(
        Red_SignaltoCheck[25]), .Z(Check1_CheckInst_0_n137) );
  XOR2_X1 Check1_CheckInst_0_U141 ( .A(Red_MC_output2[8]), .B(
        Red_SignaltoCheck[24]), .Z(Check1_CheckInst_0_n138) );
  NOR2_X1 Check1_CheckInst_0_U140 ( .A1(Check1_CheckInst_0_n136), .A2(
        Check1_CheckInst_0_n135), .ZN(Check1_CheckInst_0_n184) );
  NAND2_X1 Check1_CheckInst_0_U139 ( .A1(Check1_CheckInst_0_n134), .A2(
        Check1_CheckInst_0_n133), .ZN(Check1_CheckInst_0_n135) );
  NOR2_X1 Check1_CheckInst_0_U138 ( .A1(Check1_CheckInst_0_n132), .A2(
        Check1_CheckInst_0_n131), .ZN(Check1_CheckInst_0_n133) );
  NAND2_X1 Check1_CheckInst_0_U137 ( .A1(Check1_CheckInst_0_n130), .A2(
        Check1_CheckInst_0_n129), .ZN(Check1_CheckInst_0_n131) );
  XNOR2_X1 Check1_CheckInst_0_U136 ( .A(Red_MC_output2[11]), .B(
        Red_SignaltoCheck[27]), .ZN(Check1_CheckInst_0_n129) );
  XNOR2_X1 Check1_CheckInst_0_U135 ( .A(Red_MC_output2[7]), .B(
        Red_SignaltoCheck[23]), .ZN(Check1_CheckInst_0_n130) );
  NAND2_X1 Check1_CheckInst_0_U134 ( .A1(Check1_CheckInst_0_n128), .A2(
        Check1_CheckInst_0_n127), .ZN(Check1_CheckInst_0_n132) );
  XNOR2_X1 Check1_CheckInst_0_U133 ( .A(Red_MC_output2[10]), .B(
        Red_SignaltoCheck[26]), .ZN(Check1_CheckInst_0_n127) );
  XNOR2_X1 Check1_CheckInst_0_U132 ( .A(Red_MC_output2[12]), .B(
        Red_SignaltoCheck[28]), .ZN(Check1_CheckInst_0_n128) );
  NOR2_X1 Check1_CheckInst_0_U131 ( .A1(Check1_CheckInst_0_n126), .A2(
        Check1_CheckInst_0_n125), .ZN(Check1_CheckInst_0_n134) );
  XOR2_X1 Check1_CheckInst_0_U130 ( .A(Red_ShiftRowsOutput2[11]), .B(
        Red_SignaltoCheck[43]), .Z(Check1_CheckInst_0_n125) );
  XOR2_X1 Check1_CheckInst_0_U129 ( .A(Red_ShiftRowsOutput2[10]), .B(
        Red_SignaltoCheck[42]), .Z(Check1_CheckInst_0_n126) );
  NAND2_X1 Check1_CheckInst_0_U128 ( .A1(Check1_CheckInst_0_n124), .A2(
        Check1_CheckInst_0_n123), .ZN(Check1_CheckInst_0_n136) );
  XNOR2_X1 Check1_CheckInst_0_U127 ( .A(Red_ShiftRowsOutput2[13]), .B(
        Red_SignaltoCheck[45]), .ZN(Check1_CheckInst_0_n123) );
  XNOR2_X1 Check1_CheckInst_0_U126 ( .A(Red_ShiftRowsOutput2[9]), .B(
        Red_SignaltoCheck[41]), .ZN(Check1_CheckInst_0_n124) );
  NAND2_X1 Check1_CheckInst_0_U125 ( .A1(Check1_CheckInst_0_n122), .A2(
        Check1_CheckInst_0_n121), .ZN(Check1_CheckInst_0_n186) );
  NOR2_X1 Check1_CheckInst_0_U124 ( .A1(Check1_CheckInst_0_n120), .A2(
        Check1_CheckInst_0_n119), .ZN(Check1_CheckInst_0_n121) );
  NAND2_X1 Check1_CheckInst_0_U123 ( .A1(Check1_CheckInst_0_n118), .A2(
        Check1_CheckInst_0_n117), .ZN(Check1_CheckInst_0_n119) );
  NOR2_X1 Check1_CheckInst_0_U122 ( .A1(Check1_CheckInst_0_n116), .A2(
        Check1_CheckInst_0_n115), .ZN(Check1_CheckInst_0_n117) );
  XOR2_X1 Check1_CheckInst_0_U121 ( .A(Red_SubCellInput2[4]), .B(
        Red_SignaltoCheck[52]), .Z(Check1_CheckInst_0_n115) );
  XOR2_X1 Check1_CheckInst_0_U120 ( .A(Red_SubCellInput2[3]), .B(
        Red_SignaltoCheck[51]), .Z(Check1_CheckInst_0_n116) );
  XNOR2_X1 Check1_CheckInst_0_U119 ( .A(Red_SubCellInput2[2]), .B(
        Red_SignaltoCheck[50]), .ZN(Check1_CheckInst_0_n118) );
  NAND2_X1 Check1_CheckInst_0_U118 ( .A1(Check1_CheckInst_0_n114), .A2(
        Check1_CheckInst_0_n113), .ZN(Check1_CheckInst_0_n120) );
  NOR2_X1 Check1_CheckInst_0_U117 ( .A1(Check1_CheckInst_0_n112), .A2(
        Check1_CheckInst_0_n111), .ZN(Check1_CheckInst_0_n113) );
  NAND2_X1 Check1_CheckInst_0_U116 ( .A1(Check1_CheckInst_0_n110), .A2(
        Check1_CheckInst_0_n109), .ZN(Check1_CheckInst_0_n111) );
  NOR2_X1 Check1_CheckInst_0_U115 ( .A1(Check1_CheckInst_0_n108), .A2(
        Check1_CheckInst_0_n107), .ZN(Check1_CheckInst_0_n109) );
  XOR2_X1 Check1_CheckInst_0_U114 ( .A(Red_MC_output[2]), .B(
        Red_SignaltoCheck[66]), .Z(Check1_CheckInst_0_n107) );
  XOR2_X1 Check1_CheckInst_0_U113 ( .A(Red_MC_output[4]), .B(
        Red_SignaltoCheck[68]), .Z(Check1_CheckInst_0_n108) );
  XNOR2_X1 Check1_CheckInst_0_U112 ( .A(Red_MC_output[3]), .B(
        Red_SignaltoCheck[67]), .ZN(Check1_CheckInst_0_n110) );
  NAND2_X1 Check1_CheckInst_0_U111 ( .A1(Check1_CheckInst_0_n106), .A2(
        Check1_CheckInst_0_n105), .ZN(Check1_CheckInst_0_n112) );
  NOR2_X1 Check1_CheckInst_0_U110 ( .A1(Check1_CheckInst_0_n104), .A2(
        Check1_CheckInst_0_n103), .ZN(Check1_CheckInst_0_n105) );
  NAND2_X1 Check1_CheckInst_0_U109 ( .A1(Check1_CheckInst_0_n102), .A2(
        Check1_CheckInst_0_n101), .ZN(Check1_CheckInst_0_n103) );
  NOR2_X1 Check1_CheckInst_0_U108 ( .A1(Check1_CheckInst_0_n100), .A2(
        Check1_CheckInst_0_n99), .ZN(Check1_CheckInst_0_n101) );
  XOR2_X1 Check1_CheckInst_0_U107 ( .A(Red_SubCellInput2[11]), .B(
        Red_SignaltoCheck[59]), .Z(Check1_CheckInst_0_n99) );
  XOR2_X1 Check1_CheckInst_0_U106 ( .A(Red_SubCellInput2[13]), .B(
        Red_SignaltoCheck[61]), .Z(Check1_CheckInst_0_n100) );
  XNOR2_X1 Check1_CheckInst_0_U105 ( .A(Red_MC_output[5]), .B(
        Red_SignaltoCheck[69]), .ZN(Check1_CheckInst_0_n102) );
  NAND2_X1 Check1_CheckInst_0_U104 ( .A1(Check1_CheckInst_0_n98), .A2(
        Check1_CheckInst_0_n97), .ZN(Check1_CheckInst_0_n104) );
  NOR2_X1 Check1_CheckInst_0_U103 ( .A1(Check1_CheckInst_0_n96), .A2(
        Check1_CheckInst_0_n95), .ZN(Check1_CheckInst_0_n97) );
  XOR2_X1 Check1_CheckInst_0_U102 ( .A(Red_SubCellInput2[12]), .B(
        Red_SignaltoCheck[60]), .Z(Check1_CheckInst_0_n95) );
  XOR2_X1 Check1_CheckInst_0_U101 ( .A(Red_SubCellInput2[14]), .B(
        Red_SignaltoCheck[62]), .Z(Check1_CheckInst_0_n96) );
  NOR2_X1 Check1_CheckInst_0_U100 ( .A1(Check1_CheckInst_0_n94), .A2(
        Check1_CheckInst_0_n93), .ZN(Check1_CheckInst_0_n98) );
  XOR2_X1 Check1_CheckInst_0_U99 ( .A(Red_MC_output[0]), .B(
        Red_SignaltoCheck[64]), .Z(Check1_CheckInst_0_n93) );
  XOR2_X1 Check1_CheckInst_0_U98 ( .A(Red_SubCellInput2[15]), .B(
        Red_SignaltoCheck[63]), .Z(Check1_CheckInst_0_n94) );
  XNOR2_X1 Check1_CheckInst_0_U97 ( .A(Red_SignaltoCheck[70]), .B(
        Red_MC_output[6]), .ZN(Check1_CheckInst_0_n106) );
  XNOR2_X1 Check1_CheckInst_0_U96 ( .A(Red_SignaltoCheck[65]), .B(
        Red_MC_output[1]), .ZN(Check1_CheckInst_0_n114) );
  XNOR2_X1 Check1_CheckInst_0_U95 ( .A(Red_SignaltoCheck[48]), .B(
        Red_SubCellInput2[0]), .ZN(Check1_CheckInst_0_n122) );
  NOR2_X1 Check1_CheckInst_0_U94 ( .A1(Check1_CheckInst_0_n92), .A2(
        Check1_CheckInst_0_n91), .ZN(Check1_CheckInst_0_n188) );
  NAND2_X1 Check1_CheckInst_0_U93 ( .A1(Check1_CheckInst_0_n90), .A2(
        Check1_CheckInst_0_n89), .ZN(Check1_CheckInst_0_n91) );
  NOR2_X1 Check1_CheckInst_0_U92 ( .A1(Check1_CheckInst_0_n88), .A2(
        Check1_CheckInst_0_n87), .ZN(Check1_CheckInst_0_n89) );
  NAND2_X1 Check1_CheckInst_0_U91 ( .A1(Check1_CheckInst_0_n86), .A2(
        Check1_CheckInst_0_n85), .ZN(Check1_CheckInst_0_n87) );
  NOR2_X1 Check1_CheckInst_0_U90 ( .A1(Check1_CheckInst_0_n84), .A2(
        Check1_CheckInst_0_n83), .ZN(Check1_CheckInst_0_n85) );
  NAND2_X1 Check1_CheckInst_0_U89 ( .A1(Check1_CheckInst_0_n82), .A2(
        Check1_CheckInst_0_n81), .ZN(Check1_CheckInst_0_n83) );
  NOR2_X1 Check1_CheckInst_0_U88 ( .A1(Check1_CheckInst_0_n80), .A2(
        Check1_CheckInst_0_n79), .ZN(Check1_CheckInst_0_n81) );
  XOR2_X1 Check1_CheckInst_0_U87 ( .A(Red_ShiftRowsOutput2[12]), .B(
        Red_SignaltoCheck[44]), .Z(Check1_CheckInst_0_n79) );
  XOR2_X1 Check1_CheckInst_0_U86 ( .A(Red_ShiftRowsOutput2[14]), .B(
        Red_SignaltoCheck[46]), .Z(Check1_CheckInst_0_n80) );
  NOR2_X1 Check1_CheckInst_0_U85 ( .A1(Check1_CheckInst_0_n78), .A2(
        Check1_CheckInst_0_n77), .ZN(Check1_CheckInst_0_n82) );
  XOR2_X1 Check1_CheckInst_0_U84 ( .A(Red_ShiftRowsOutput2[5]), .B(
        Red_SignaltoCheck[37]), .Z(Check1_CheckInst_0_n77) );
  XOR2_X1 Check1_CheckInst_0_U83 ( .A(Red_ShiftRowsOutput2[4]), .B(
        Red_SignaltoCheck[36]), .Z(Check1_CheckInst_0_n78) );
  NAND2_X1 Check1_CheckInst_0_U82 ( .A1(Check1_CheckInst_0_n76), .A2(
        Check1_CheckInst_0_n75), .ZN(Check1_CheckInst_0_n84) );
  XNOR2_X1 Check1_CheckInst_0_U81 ( .A(Red_ShiftRowsOutput2[7]), .B(
        Red_SignaltoCheck[39]), .ZN(Check1_CheckInst_0_n75) );
  XNOR2_X1 Check1_CheckInst_0_U80 ( .A(Red_ShiftRowsOutput2[3]), .B(
        Red_SignaltoCheck[35]), .ZN(Check1_CheckInst_0_n76) );
  NOR2_X1 Check1_CheckInst_0_U79 ( .A1(Check1_CheckInst_0_n74), .A2(
        Check1_CheckInst_0_n73), .ZN(Check1_CheckInst_0_n86) );
  XOR2_X1 Check1_CheckInst_0_U78 ( .A(Red_ShiftRowsOutput2[6]), .B(
        Red_SignaltoCheck[38]), .Z(Check1_CheckInst_0_n73) );
  XOR2_X1 Check1_CheckInst_0_U77 ( .A(Red_ShiftRowsOutput2[8]), .B(
        Red_SignaltoCheck[40]), .Z(Check1_CheckInst_0_n74) );
  NAND2_X1 Check1_CheckInst_0_U76 ( .A1(Check1_CheckInst_0_n72), .A2(
        Check1_CheckInst_0_n71), .ZN(Check1_CheckInst_0_n88) );
  NOR2_X1 Check1_CheckInst_0_U75 ( .A1(Check1_CheckInst_0_n70), .A2(
        Check1_CheckInst_0_n69), .ZN(Check1_CheckInst_0_n71) );
  NAND2_X1 Check1_CheckInst_0_U74 ( .A1(Check1_CheckInst_0_n68), .A2(
        Check1_CheckInst_0_n67), .ZN(Check1_CheckInst_0_n69) );
  NOR2_X1 Check1_CheckInst_0_U73 ( .A1(Check1_CheckInst_0_n66), .A2(
        Check1_CheckInst_0_n65), .ZN(Check1_CheckInst_0_n67) );
  XOR2_X1 Check1_CheckInst_0_U72 ( .A(Red_AddRoundKeyOutput[7]), .B(
        Red_SignaltoCheck[7]), .Z(Check1_CheckInst_0_n65) );
  XOR2_X1 Check1_CheckInst_0_U71 ( .A(Red_AddRoundKeyOutput[6]), .B(
        Red_SignaltoCheck[6]), .Z(Check1_CheckInst_0_n66) );
  NOR2_X1 Check1_CheckInst_0_U70 ( .A1(Check1_CheckInst_0_n64), .A2(
        Check1_CheckInst_0_n63), .ZN(Check1_CheckInst_0_n68) );
  XOR2_X1 Check1_CheckInst_0_U69 ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[9]), .Z(Check1_CheckInst_0_n63) );
  XOR2_X1 Check1_CheckInst_0_U68 ( .A(Red_AddRoundKeyOutput[5]), .B(
        Red_SignaltoCheck[5]), .Z(Check1_CheckInst_0_n64) );
  NAND2_X1 Check1_CheckInst_0_U67 ( .A1(Check1_CheckInst_0_n62), .A2(
        Check1_CheckInst_0_n61), .ZN(Check1_CheckInst_0_n70) );
  XNOR2_X1 Check1_CheckInst_0_U66 ( .A(Red_AddRoundKeyOutput[8]), .B(
        Red_SignaltoCheck[8]), .ZN(Check1_CheckInst_0_n61) );
  XNOR2_X1 Check1_CheckInst_0_U65 ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[10]), .ZN(Check1_CheckInst_0_n62) );
  NOR2_X1 Check1_CheckInst_0_U64 ( .A1(Check1_CheckInst_0_n60), .A2(
        Check1_CheckInst_0_n59), .ZN(Check1_CheckInst_0_n72) );
  XOR2_X1 Check1_CheckInst_0_U63 ( .A(Red_ShiftRowsOutput[15]), .B(
        Red_SignaltoCheck[95]), .Z(Check1_CheckInst_0_n59) );
  XOR2_X1 Check1_CheckInst_0_U62 ( .A(Red_SignaltoCheck[1]), .B(
        Red_AddRoundKeyOutput[1]), .Z(Check1_CheckInst_0_n60) );
  NOR2_X1 Check1_CheckInst_0_U61 ( .A1(Check1_CheckInst_0_n58), .A2(
        Check1_CheckInst_0_n57), .ZN(Check1_CheckInst_0_n90) );
  NAND2_X1 Check1_CheckInst_0_U60 ( .A1(Check1_CheckInst_0_n56), .A2(
        Check1_CheckInst_0_n55), .ZN(Check1_CheckInst_0_n57) );
  NOR2_X1 Check1_CheckInst_0_U59 ( .A1(Check1_CheckInst_0_n54), .A2(
        Check1_CheckInst_0_n53), .ZN(Check1_CheckInst_0_n55) );
  NAND2_X1 Check1_CheckInst_0_U58 ( .A1(Check1_CheckInst_0_n52), .A2(
        Check1_CheckInst_0_n51), .ZN(Check1_CheckInst_0_n53) );
  XNOR2_X1 Check1_CheckInst_0_U57 ( .A(Red_AddRoundKeyOutput[3]), .B(
        Red_SignaltoCheck[3]), .ZN(Check1_CheckInst_0_n51) );
  XNOR2_X1 Check1_CheckInst_0_U56 ( .A(Red_SignaltoCheck[0]), .B(
        Red_AddRoundKeyOutput[0]), .ZN(Check1_CheckInst_0_n52) );
  NAND2_X1 Check1_CheckInst_0_U55 ( .A1(Check1_CheckInst_0_n50), .A2(
        Check1_CheckInst_0_n49), .ZN(Check1_CheckInst_0_n54) );
  XNOR2_X1 Check1_CheckInst_0_U54 ( .A(Red_AddRoundKeyOutput[2]), .B(
        Red_SignaltoCheck[2]), .ZN(Check1_CheckInst_0_n49) );
  XNOR2_X1 Check1_CheckInst_0_U53 ( .A(Red_AddRoundKeyOutput[4]), .B(
        Red_SignaltoCheck[4]), .ZN(Check1_CheckInst_0_n50) );
  NOR2_X1 Check1_CheckInst_0_U52 ( .A1(Check1_CheckInst_0_n48), .A2(
        Check1_CheckInst_0_n47), .ZN(Check1_CheckInst_0_n56) );
  XOR2_X1 Check1_CheckInst_0_U51 ( .A(Red_MC_output2[3]), .B(
        Red_SignaltoCheck[19]), .Z(Check1_CheckInst_0_n47) );
  XOR2_X1 Check1_CheckInst_0_U50 ( .A(Red_MC_output2[2]), .B(
        Red_SignaltoCheck[18]), .Z(Check1_CheckInst_0_n48) );
  NAND2_X1 Check1_CheckInst_0_U49 ( .A1(Check1_CheckInst_0_n46), .A2(
        Check1_CheckInst_0_n45), .ZN(Check1_CheckInst_0_n58) );
  XNOR2_X1 Check1_CheckInst_0_U48 ( .A(Red_MC_output2[5]), .B(
        Red_SignaltoCheck[21]), .ZN(Check1_CheckInst_0_n45) );
  XNOR2_X1 Check1_CheckInst_0_U47 ( .A(Red_MC_output2[1]), .B(
        Red_SignaltoCheck[17]), .ZN(Check1_CheckInst_0_n46) );
  NAND2_X1 Check1_CheckInst_0_U46 ( .A1(Check1_CheckInst_0_n44), .A2(
        Check1_CheckInst_0_n43), .ZN(Check1_CheckInst_0_n92) );
  NOR2_X1 Check1_CheckInst_0_U45 ( .A1(Check1_CheckInst_0_n42), .A2(
        Check1_CheckInst_0_n41), .ZN(Check1_CheckInst_0_n43) );
  NAND2_X1 Check1_CheckInst_0_U44 ( .A1(Check1_CheckInst_0_n40), .A2(
        Check1_CheckInst_0_n39), .ZN(Check1_CheckInst_0_n41) );
  NOR2_X1 Check1_CheckInst_0_U43 ( .A1(Check1_CheckInst_0_n38), .A2(
        Check1_CheckInst_0_n37), .ZN(Check1_CheckInst_0_n39) );
  XOR2_X1 Check1_CheckInst_0_U42 ( .A(Red_MC_output2[4]), .B(
        Red_SignaltoCheck[20]), .Z(Check1_CheckInst_0_n37) );
  XOR2_X1 Check1_CheckInst_0_U41 ( .A(Red_MC_output2[6]), .B(
        Red_SignaltoCheck[22]), .Z(Check1_CheckInst_0_n38) );
  NOR2_X1 Check1_CheckInst_0_U40 ( .A1(Check1_CheckInst_0_n36), .A2(
        Check1_CheckInst_0_n35), .ZN(Check1_CheckInst_0_n40) );
  XOR2_X1 Check1_CheckInst_0_U39 ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[13]), .Z(Check1_CheckInst_0_n35) );
  XOR2_X1 Check1_CheckInst_0_U38 ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[12]), .Z(Check1_CheckInst_0_n36) );
  NAND2_X1 Check1_CheckInst_0_U37 ( .A1(Check1_CheckInst_0_n34), .A2(
        Check1_CheckInst_0_n33), .ZN(Check1_CheckInst_0_n42) );
  XNOR2_X1 Check1_CheckInst_0_U36 ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[15]), .ZN(Check1_CheckInst_0_n33) );
  XNOR2_X1 Check1_CheckInst_0_U35 ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[11]), .ZN(Check1_CheckInst_0_n34) );
  NOR2_X1 Check1_CheckInst_0_U34 ( .A1(Check1_CheckInst_0_n32), .A2(
        Check1_CheckInst_0_n31), .ZN(Check1_CheckInst_0_n44) );
  XOR2_X1 Check1_CheckInst_0_U33 ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[14]), .Z(Check1_CheckInst_0_n31) );
  XOR2_X1 Check1_CheckInst_0_U32 ( .A(Red_MC_output2[0]), .B(
        Red_SignaltoCheck[16]), .Z(Check1_CheckInst_0_n32) );
  NAND2_X1 Check1_CheckInst_0_U31 ( .A1(Check1_CheckInst_0_n30), .A2(
        Check1_CheckInst_0_n29), .ZN(Check1_CheckInst_0_n190) );
  NOR2_X1 Check1_CheckInst_0_U30 ( .A1(Check1_CheckInst_0_n28), .A2(
        Check1_CheckInst_0_n27), .ZN(Check1_CheckInst_0_n29) );
  NAND2_X1 Check1_CheckInst_0_U29 ( .A1(Check1_CheckInst_0_n26), .A2(
        Check1_CheckInst_0_n25), .ZN(Check1_CheckInst_0_n27) );
  NOR2_X1 Check1_CheckInst_0_U28 ( .A1(Check1_CheckInst_0_n24), .A2(
        Check1_CheckInst_0_n23), .ZN(Check1_CheckInst_0_n25) );
  XOR2_X1 Check1_CheckInst_0_U27 ( .A(Red_ShiftRowsOutput[3]), .B(
        Red_SignaltoCheck[83]), .Z(Check1_CheckInst_0_n23) );
  XOR2_X1 Check1_CheckInst_0_U26 ( .A(Red_ShiftRowsOutput[5]), .B(
        Red_SignaltoCheck[85]), .Z(Check1_CheckInst_0_n24) );
  XNOR2_X1 Check1_CheckInst_0_U25 ( .A(Red_ShiftRowsOutput[13]), .B(
        Red_SignaltoCheck[93]), .ZN(Check1_CheckInst_0_n26) );
  NAND2_X1 Check1_CheckInst_0_U24 ( .A1(Check1_CheckInst_0_n22), .A2(
        Check1_CheckInst_0_n21), .ZN(Check1_CheckInst_0_n28) );
  NOR2_X1 Check1_CheckInst_0_U23 ( .A1(Check1_CheckInst_0_n20), .A2(
        Check1_CheckInst_0_n19), .ZN(Check1_CheckInst_0_n21) );
  NAND2_X1 Check1_CheckInst_0_U22 ( .A1(Check1_CheckInst_0_n18), .A2(
        Check1_CheckInst_0_n17), .ZN(Check1_CheckInst_0_n19) );
  NOR2_X1 Check1_CheckInst_0_U21 ( .A1(Check1_CheckInst_0_n16), .A2(
        Check1_CheckInst_0_n15), .ZN(Check1_CheckInst_0_n17) );
  XOR2_X1 Check1_CheckInst_0_U20 ( .A(Red_ShiftRowsOutput[8]), .B(
        Red_SignaltoCheck[88]), .Z(Check1_CheckInst_0_n15) );
  XOR2_X1 Check1_CheckInst_0_U19 ( .A(Red_ShiftRowsOutput[7]), .B(
        Red_SignaltoCheck[87]), .Z(Check1_CheckInst_0_n16) );
  XNOR2_X1 Check1_CheckInst_0_U18 ( .A(Red_ShiftRowsOutput[6]), .B(
        Red_SignaltoCheck[86]), .ZN(Check1_CheckInst_0_n18) );
  NAND2_X1 Check1_CheckInst_0_U17 ( .A1(Check1_CheckInst_0_n14), .A2(
        Check1_CheckInst_0_n13), .ZN(Check1_CheckInst_0_n20) );
  NOR2_X1 Check1_CheckInst_0_U16 ( .A1(Check1_CheckInst_0_n12), .A2(
        Check1_CheckInst_0_n11), .ZN(Check1_CheckInst_0_n13) );
  NAND2_X1 Check1_CheckInst_0_U15 ( .A1(Check1_CheckInst_0_n10), .A2(
        Check1_CheckInst_0_n9), .ZN(Check1_CheckInst_0_n11) );
  NOR2_X1 Check1_CheckInst_0_U14 ( .A1(Check1_CheckInst_0_n8), .A2(
        Check1_CheckInst_0_n7), .ZN(Check1_CheckInst_0_n9) );
  XOR2_X1 Check1_CheckInst_0_U13 ( .A(Red_SubCellInput2[6]), .B(
        Red_SignaltoCheck[54]), .Z(Check1_CheckInst_0_n7) );
  XOR2_X1 Check1_CheckInst_0_U12 ( .A(Red_SubCellInput2[8]), .B(
        Red_SignaltoCheck[56]), .Z(Check1_CheckInst_0_n8) );
  XNOR2_X1 Check1_CheckInst_0_U11 ( .A(Red_SubCellInput2[7]), .B(
        Red_SignaltoCheck[55]), .ZN(Check1_CheckInst_0_n10) );
  NAND2_X1 Check1_CheckInst_0_U10 ( .A1(Check1_CheckInst_0_n6), .A2(
        Check1_CheckInst_0_n5), .ZN(Check1_CheckInst_0_n12) );
  NOR2_X1 Check1_CheckInst_0_U9 ( .A1(Check1_CheckInst_0_n4), .A2(
        Check1_CheckInst_0_n3), .ZN(Check1_CheckInst_0_n5) );
  XOR2_X1 Check1_CheckInst_0_U8 ( .A(Red_SubCellInput2[10]), .B(
        Red_SignaltoCheck[58]), .Z(Check1_CheckInst_0_n3) );
  XOR2_X1 Check1_CheckInst_0_U7 ( .A(Red_SubCellInput2[9]), .B(
        Red_SignaltoCheck[57]), .Z(Check1_CheckInst_0_n4) );
  NOR2_X1 Check1_CheckInst_0_U6 ( .A1(Check1_CheckInst_0_n2), .A2(
        Check1_CheckInst_0_n1), .ZN(Check1_CheckInst_0_n6) );
  XOR2_X1 Check1_CheckInst_0_U5 ( .A(Red_ShiftRowsOutput2[15]), .B(
        Red_SignaltoCheck[47]), .Z(Check1_CheckInst_0_n1) );
  XOR2_X1 Check1_CheckInst_0_U4 ( .A(Red_SubCellInput2[1]), .B(
        Red_SignaltoCheck[49]), .Z(Check1_CheckInst_0_n2) );
  XNOR2_X1 Check1_CheckInst_0_U3 ( .A(Red_SignaltoCheck[53]), .B(
        Red_SubCellInput2[5]), .ZN(Check1_CheckInst_0_n14) );
  XNOR2_X1 Check1_CheckInst_0_U2 ( .A(Red_SignaltoCheck[84]), .B(
        Red_ShiftRowsOutput[4]), .ZN(Check1_CheckInst_0_n22) );
  XNOR2_X1 Check1_CheckInst_0_U1 ( .A(Red_SignaltoCheck[94]), .B(
        Red_ShiftRowsOutput[14]), .ZN(Check1_CheckInst_0_n30) );
endmodule

