
module LED64Enc ( clk, Plaintext, Key, Ciphertext, ErrorFlag );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* fiver="clock" *)input clk;
  output ErrorFlag;
  wire   n4, SubCellInst_LFInst_0_LFInst_0_n9,
         SubCellInst_LFInst_0_LFInst_0_n8, SubCellInst_LFInst_0_LFInst_0_n7,
         SubCellInst_LFInst_0_LFInst_0_n10, SubCellInst_LFInst_0_LFInst_1_n26,
         SubCellInst_LFInst_0_LFInst_1_n25, SubCellInst_LFInst_0_LFInst_1_n24,
         SubCellInst_LFInst_0_LFInst_1_n23, SubCellInst_LFInst_0_LFInst_1_n22,
         SubCellInst_LFInst_0_LFInst_1_n21, SubCellInst_LFInst_0_LFInst_1_n20,
         SubCellInst_LFInst_0_LFInst_1_n19, SubCellInst_LFInst_0_LFInst_1_n18,
         SubCellInst_LFInst_0_LFInst_2_n28, SubCellInst_LFInst_0_LFInst_2_n27,
         SubCellInst_LFInst_0_LFInst_2_n26, SubCellInst_LFInst_0_LFInst_2_n25,
         SubCellInst_LFInst_0_LFInst_2_n24, SubCellInst_LFInst_0_LFInst_2_n23,
         SubCellInst_LFInst_0_LFInst_2_n22, SubCellInst_LFInst_0_LFInst_3_n26,
         SubCellInst_LFInst_0_LFInst_3_n25, SubCellInst_LFInst_0_LFInst_3_n24,
         SubCellInst_LFInst_0_LFInst_3_n23, SubCellInst_LFInst_0_LFInst_3_n22,
         SubCellInst_LFInst_0_LFInst_3_n21, SubCellInst_LFInst_0_LFInst_3_n20,
         SubCellInst_LFInst_0_LFInst_3_n19, SubCellInst_LFInst_1_LFInst_0_n9,
         SubCellInst_LFInst_1_LFInst_0_n8, SubCellInst_LFInst_1_LFInst_0_n7,
         SubCellInst_LFInst_1_LFInst_0_n10, SubCellInst_LFInst_1_LFInst_1_n26,
         SubCellInst_LFInst_1_LFInst_1_n25, SubCellInst_LFInst_1_LFInst_1_n24,
         SubCellInst_LFInst_1_LFInst_1_n23, SubCellInst_LFInst_1_LFInst_1_n22,
         SubCellInst_LFInst_1_LFInst_1_n21, SubCellInst_LFInst_1_LFInst_1_n20,
         SubCellInst_LFInst_1_LFInst_1_n19, SubCellInst_LFInst_1_LFInst_1_n18,
         SubCellInst_LFInst_1_LFInst_2_n28, SubCellInst_LFInst_1_LFInst_2_n27,
         SubCellInst_LFInst_1_LFInst_2_n26, SubCellInst_LFInst_1_LFInst_2_n25,
         SubCellInst_LFInst_1_LFInst_2_n24, SubCellInst_LFInst_1_LFInst_2_n23,
         SubCellInst_LFInst_1_LFInst_2_n22, SubCellInst_LFInst_1_LFInst_3_n26,
         SubCellInst_LFInst_1_LFInst_3_n25, SubCellInst_LFInst_1_LFInst_3_n24,
         SubCellInst_LFInst_1_LFInst_3_n23, SubCellInst_LFInst_1_LFInst_3_n22,
         SubCellInst_LFInst_1_LFInst_3_n21, SubCellInst_LFInst_1_LFInst_3_n20,
         SubCellInst_LFInst_1_LFInst_3_n19, SubCellInst_LFInst_2_LFInst_0_n9,
         SubCellInst_LFInst_2_LFInst_0_n8, SubCellInst_LFInst_2_LFInst_0_n7,
         SubCellInst_LFInst_2_LFInst_0_n10, SubCellInst_LFInst_2_LFInst_1_n26,
         SubCellInst_LFInst_2_LFInst_1_n25, SubCellInst_LFInst_2_LFInst_1_n24,
         SubCellInst_LFInst_2_LFInst_1_n23, SubCellInst_LFInst_2_LFInst_1_n22,
         SubCellInst_LFInst_2_LFInst_1_n21, SubCellInst_LFInst_2_LFInst_1_n20,
         SubCellInst_LFInst_2_LFInst_1_n19, SubCellInst_LFInst_2_LFInst_1_n18,
         SubCellInst_LFInst_2_LFInst_2_n28, SubCellInst_LFInst_2_LFInst_2_n27,
         SubCellInst_LFInst_2_LFInst_2_n26, SubCellInst_LFInst_2_LFInst_2_n25,
         SubCellInst_LFInst_2_LFInst_2_n24, SubCellInst_LFInst_2_LFInst_2_n23,
         SubCellInst_LFInst_2_LFInst_2_n22, SubCellInst_LFInst_2_LFInst_3_n26,
         SubCellInst_LFInst_2_LFInst_3_n25, SubCellInst_LFInst_2_LFInst_3_n24,
         SubCellInst_LFInst_2_LFInst_3_n23, SubCellInst_LFInst_2_LFInst_3_n22,
         SubCellInst_LFInst_2_LFInst_3_n21, SubCellInst_LFInst_2_LFInst_3_n20,
         SubCellInst_LFInst_2_LFInst_3_n19, SubCellInst_LFInst_3_LFInst_0_n9,
         SubCellInst_LFInst_3_LFInst_0_n8, SubCellInst_LFInst_3_LFInst_0_n7,
         SubCellInst_LFInst_3_LFInst_0_n10, SubCellInst_LFInst_3_LFInst_1_n26,
         SubCellInst_LFInst_3_LFInst_1_n25, SubCellInst_LFInst_3_LFInst_1_n24,
         SubCellInst_LFInst_3_LFInst_1_n23, SubCellInst_LFInst_3_LFInst_1_n22,
         SubCellInst_LFInst_3_LFInst_1_n21, SubCellInst_LFInst_3_LFInst_1_n20,
         SubCellInst_LFInst_3_LFInst_1_n19, SubCellInst_LFInst_3_LFInst_1_n18,
         SubCellInst_LFInst_3_LFInst_2_n28, SubCellInst_LFInst_3_LFInst_2_n27,
         SubCellInst_LFInst_3_LFInst_2_n26, SubCellInst_LFInst_3_LFInst_2_n25,
         SubCellInst_LFInst_3_LFInst_2_n24, SubCellInst_LFInst_3_LFInst_2_n23,
         SubCellInst_LFInst_3_LFInst_2_n22, SubCellInst_LFInst_3_LFInst_3_n26,
         SubCellInst_LFInst_3_LFInst_3_n25, SubCellInst_LFInst_3_LFInst_3_n24,
         SubCellInst_LFInst_3_LFInst_3_n23, SubCellInst_LFInst_3_LFInst_3_n22,
         SubCellInst_LFInst_3_LFInst_3_n21, SubCellInst_LFInst_3_LFInst_3_n20,
         SubCellInst_LFInst_3_LFInst_3_n19, SubCellInst_LFInst_4_LFInst_0_n8,
         SubCellInst_LFInst_4_LFInst_0_n7, SubCellInst_LFInst_4_LFInst_0_n6,
         SubCellInst_LFInst_4_LFInst_1_n26, SubCellInst_LFInst_4_LFInst_1_n25,
         SubCellInst_LFInst_4_LFInst_1_n24, SubCellInst_LFInst_4_LFInst_1_n23,
         SubCellInst_LFInst_4_LFInst_1_n22, SubCellInst_LFInst_4_LFInst_1_n21,
         SubCellInst_LFInst_4_LFInst_1_n20, SubCellInst_LFInst_4_LFInst_1_n19,
         SubCellInst_LFInst_4_LFInst_1_n18, SubCellInst_LFInst_4_LFInst_2_n29,
         SubCellInst_LFInst_4_LFInst_2_n28, SubCellInst_LFInst_4_LFInst_2_n27,
         SubCellInst_LFInst_4_LFInst_2_n26, SubCellInst_LFInst_4_LFInst_2_n25,
         SubCellInst_LFInst_4_LFInst_2_n24, SubCellInst_LFInst_4_LFInst_2_n23,
         SubCellInst_LFInst_4_LFInst_2_n22, SubCellInst_LFInst_4_LFInst_3_n26,
         SubCellInst_LFInst_4_LFInst_3_n25, SubCellInst_LFInst_4_LFInst_3_n24,
         SubCellInst_LFInst_4_LFInst_3_n23, SubCellInst_LFInst_4_LFInst_3_n22,
         SubCellInst_LFInst_4_LFInst_3_n21, SubCellInst_LFInst_4_LFInst_3_n20,
         SubCellInst_LFInst_4_LFInst_3_n19, SubCellInst_LFInst_5_LFInst_0_n8,
         SubCellInst_LFInst_5_LFInst_0_n7, SubCellInst_LFInst_5_LFInst_0_n6,
         SubCellInst_LFInst_5_LFInst_1_n26, SubCellInst_LFInst_5_LFInst_1_n25,
         SubCellInst_LFInst_5_LFInst_1_n24, SubCellInst_LFInst_5_LFInst_1_n23,
         SubCellInst_LFInst_5_LFInst_1_n22, SubCellInst_LFInst_5_LFInst_1_n21,
         SubCellInst_LFInst_5_LFInst_1_n20, SubCellInst_LFInst_5_LFInst_1_n19,
         SubCellInst_LFInst_5_LFInst_1_n18, SubCellInst_LFInst_5_LFInst_2_n29,
         SubCellInst_LFInst_5_LFInst_2_n28, SubCellInst_LFInst_5_LFInst_2_n27,
         SubCellInst_LFInst_5_LFInst_2_n26, SubCellInst_LFInst_5_LFInst_2_n25,
         SubCellInst_LFInst_5_LFInst_2_n24, SubCellInst_LFInst_5_LFInst_2_n23,
         SubCellInst_LFInst_5_LFInst_2_n22, SubCellInst_LFInst_5_LFInst_3_n26,
         SubCellInst_LFInst_5_LFInst_3_n25, SubCellInst_LFInst_5_LFInst_3_n24,
         SubCellInst_LFInst_5_LFInst_3_n23, SubCellInst_LFInst_5_LFInst_3_n22,
         SubCellInst_LFInst_5_LFInst_3_n21, SubCellInst_LFInst_5_LFInst_3_n20,
         SubCellInst_LFInst_5_LFInst_3_n19, SubCellInst_LFInst_6_LFInst_0_n8,
         SubCellInst_LFInst_6_LFInst_0_n7, SubCellInst_LFInst_6_LFInst_0_n6,
         SubCellInst_LFInst_6_LFInst_1_n26, SubCellInst_LFInst_6_LFInst_1_n25,
         SubCellInst_LFInst_6_LFInst_1_n24, SubCellInst_LFInst_6_LFInst_1_n23,
         SubCellInst_LFInst_6_LFInst_1_n22, SubCellInst_LFInst_6_LFInst_1_n21,
         SubCellInst_LFInst_6_LFInst_1_n20, SubCellInst_LFInst_6_LFInst_1_n19,
         SubCellInst_LFInst_6_LFInst_1_n18, SubCellInst_LFInst_6_LFInst_2_n29,
         SubCellInst_LFInst_6_LFInst_2_n28, SubCellInst_LFInst_6_LFInst_2_n27,
         SubCellInst_LFInst_6_LFInst_2_n26, SubCellInst_LFInst_6_LFInst_2_n25,
         SubCellInst_LFInst_6_LFInst_2_n24, SubCellInst_LFInst_6_LFInst_2_n23,
         SubCellInst_LFInst_6_LFInst_2_n22, SubCellInst_LFInst_6_LFInst_3_n26,
         SubCellInst_LFInst_6_LFInst_3_n25, SubCellInst_LFInst_6_LFInst_3_n24,
         SubCellInst_LFInst_6_LFInst_3_n23, SubCellInst_LFInst_6_LFInst_3_n22,
         SubCellInst_LFInst_6_LFInst_3_n21, SubCellInst_LFInst_6_LFInst_3_n20,
         SubCellInst_LFInst_6_LFInst_3_n19, SubCellInst_LFInst_7_LFInst_0_n8,
         SubCellInst_LFInst_7_LFInst_0_n7, SubCellInst_LFInst_7_LFInst_0_n6,
         SubCellInst_LFInst_7_LFInst_1_n26, SubCellInst_LFInst_7_LFInst_1_n25,
         SubCellInst_LFInst_7_LFInst_1_n24, SubCellInst_LFInst_7_LFInst_1_n23,
         SubCellInst_LFInst_7_LFInst_1_n22, SubCellInst_LFInst_7_LFInst_1_n21,
         SubCellInst_LFInst_7_LFInst_1_n20, SubCellInst_LFInst_7_LFInst_1_n19,
         SubCellInst_LFInst_7_LFInst_1_n18, SubCellInst_LFInst_7_LFInst_2_n29,
         SubCellInst_LFInst_7_LFInst_2_n28, SubCellInst_LFInst_7_LFInst_2_n27,
         SubCellInst_LFInst_7_LFInst_2_n26, SubCellInst_LFInst_7_LFInst_2_n25,
         SubCellInst_LFInst_7_LFInst_2_n24, SubCellInst_LFInst_7_LFInst_2_n23,
         SubCellInst_LFInst_7_LFInst_2_n22, SubCellInst_LFInst_7_LFInst_3_n26,
         SubCellInst_LFInst_7_LFInst_3_n25, SubCellInst_LFInst_7_LFInst_3_n24,
         SubCellInst_LFInst_7_LFInst_3_n23, SubCellInst_LFInst_7_LFInst_3_n22,
         SubCellInst_LFInst_7_LFInst_3_n21, SubCellInst_LFInst_7_LFInst_3_n20,
         SubCellInst_LFInst_7_LFInst_3_n19, SubCellInst_LFInst_8_LFInst_0_n11,
         SubCellInst_LFInst_8_LFInst_0_n10, SubCellInst_LFInst_8_LFInst_0_n9,
         SubCellInst_LFInst_8_LFInst_0_n12, SubCellInst_LFInst_8_LFInst_1_n26,
         SubCellInst_LFInst_8_LFInst_1_n25, SubCellInst_LFInst_8_LFInst_1_n24,
         SubCellInst_LFInst_8_LFInst_1_n23, SubCellInst_LFInst_8_LFInst_1_n22,
         SubCellInst_LFInst_8_LFInst_1_n21, SubCellInst_LFInst_8_LFInst_1_n20,
         SubCellInst_LFInst_8_LFInst_1_n19, SubCellInst_LFInst_8_LFInst_1_n18,
         SubCellInst_LFInst_8_LFInst_2_n28, SubCellInst_LFInst_8_LFInst_2_n27,
         SubCellInst_LFInst_8_LFInst_2_n26, SubCellInst_LFInst_8_LFInst_2_n25,
         SubCellInst_LFInst_8_LFInst_2_n24, SubCellInst_LFInst_8_LFInst_2_n23,
         SubCellInst_LFInst_8_LFInst_2_n22, SubCellInst_LFInst_8_LFInst_3_n26,
         SubCellInst_LFInst_8_LFInst_3_n25, SubCellInst_LFInst_8_LFInst_3_n24,
         SubCellInst_LFInst_8_LFInst_3_n23, SubCellInst_LFInst_8_LFInst_3_n22,
         SubCellInst_LFInst_8_LFInst_3_n21, SubCellInst_LFInst_8_LFInst_3_n20,
         SubCellInst_LFInst_8_LFInst_3_n19, SubCellInst_LFInst_9_LFInst_0_n12,
         SubCellInst_LFInst_9_LFInst_0_n11, SubCellInst_LFInst_9_LFInst_0_n10,
         SubCellInst_LFInst_9_LFInst_0_n9, SubCellInst_LFInst_9_LFInst_1_n26,
         SubCellInst_LFInst_9_LFInst_1_n25, SubCellInst_LFInst_9_LFInst_1_n24,
         SubCellInst_LFInst_9_LFInst_1_n23, SubCellInst_LFInst_9_LFInst_1_n22,
         SubCellInst_LFInst_9_LFInst_1_n21, SubCellInst_LFInst_9_LFInst_1_n20,
         SubCellInst_LFInst_9_LFInst_1_n19, SubCellInst_LFInst_9_LFInst_1_n18,
         SubCellInst_LFInst_9_LFInst_2_n28, SubCellInst_LFInst_9_LFInst_2_n27,
         SubCellInst_LFInst_9_LFInst_2_n26, SubCellInst_LFInst_9_LFInst_2_n25,
         SubCellInst_LFInst_9_LFInst_2_n24, SubCellInst_LFInst_9_LFInst_2_n23,
         SubCellInst_LFInst_9_LFInst_2_n22, SubCellInst_LFInst_9_LFInst_3_n26,
         SubCellInst_LFInst_9_LFInst_3_n25, SubCellInst_LFInst_9_LFInst_3_n24,
         SubCellInst_LFInst_9_LFInst_3_n23, SubCellInst_LFInst_9_LFInst_3_n22,
         SubCellInst_LFInst_9_LFInst_3_n21, SubCellInst_LFInst_9_LFInst_3_n20,
         SubCellInst_LFInst_9_LFInst_3_n19, SubCellInst_LFInst_10_LFInst_0_n12,
         SubCellInst_LFInst_10_LFInst_0_n11,
         SubCellInst_LFInst_10_LFInst_0_n10, SubCellInst_LFInst_10_LFInst_0_n9,
         SubCellInst_LFInst_10_LFInst_1_n26,
         SubCellInst_LFInst_10_LFInst_1_n25,
         SubCellInst_LFInst_10_LFInst_1_n24,
         SubCellInst_LFInst_10_LFInst_1_n23,
         SubCellInst_LFInst_10_LFInst_1_n22,
         SubCellInst_LFInst_10_LFInst_1_n21,
         SubCellInst_LFInst_10_LFInst_1_n20,
         SubCellInst_LFInst_10_LFInst_1_n19,
         SubCellInst_LFInst_10_LFInst_1_n18,
         SubCellInst_LFInst_10_LFInst_2_n28,
         SubCellInst_LFInst_10_LFInst_2_n27,
         SubCellInst_LFInst_10_LFInst_2_n26,
         SubCellInst_LFInst_10_LFInst_2_n25,
         SubCellInst_LFInst_10_LFInst_2_n24,
         SubCellInst_LFInst_10_LFInst_2_n23,
         SubCellInst_LFInst_10_LFInst_2_n22,
         SubCellInst_LFInst_10_LFInst_3_n26,
         SubCellInst_LFInst_10_LFInst_3_n25,
         SubCellInst_LFInst_10_LFInst_3_n24,
         SubCellInst_LFInst_10_LFInst_3_n23,
         SubCellInst_LFInst_10_LFInst_3_n22,
         SubCellInst_LFInst_10_LFInst_3_n21,
         SubCellInst_LFInst_10_LFInst_3_n20,
         SubCellInst_LFInst_10_LFInst_3_n19,
         SubCellInst_LFInst_11_LFInst_0_n12,
         SubCellInst_LFInst_11_LFInst_0_n11,
         SubCellInst_LFInst_11_LFInst_0_n10, SubCellInst_LFInst_11_LFInst_0_n9,
         SubCellInst_LFInst_11_LFInst_1_n26,
         SubCellInst_LFInst_11_LFInst_1_n25,
         SubCellInst_LFInst_11_LFInst_1_n24,
         SubCellInst_LFInst_11_LFInst_1_n23,
         SubCellInst_LFInst_11_LFInst_1_n22,
         SubCellInst_LFInst_11_LFInst_1_n21,
         SubCellInst_LFInst_11_LFInst_1_n20,
         SubCellInst_LFInst_11_LFInst_1_n19,
         SubCellInst_LFInst_11_LFInst_1_n18,
         SubCellInst_LFInst_11_LFInst_2_n28,
         SubCellInst_LFInst_11_LFInst_2_n27,
         SubCellInst_LFInst_11_LFInst_2_n26,
         SubCellInst_LFInst_11_LFInst_2_n25,
         SubCellInst_LFInst_11_LFInst_2_n24,
         SubCellInst_LFInst_11_LFInst_2_n23,
         SubCellInst_LFInst_11_LFInst_2_n22,
         SubCellInst_LFInst_11_LFInst_3_n26,
         SubCellInst_LFInst_11_LFInst_3_n25,
         SubCellInst_LFInst_11_LFInst_3_n24,
         SubCellInst_LFInst_11_LFInst_3_n23,
         SubCellInst_LFInst_11_LFInst_3_n22,
         SubCellInst_LFInst_11_LFInst_3_n21,
         SubCellInst_LFInst_11_LFInst_3_n20,
         SubCellInst_LFInst_11_LFInst_3_n19, SubCellInst_LFInst_12_LFInst_0_n8,
         SubCellInst_LFInst_12_LFInst_0_n7, SubCellInst_LFInst_12_LFInst_0_n6,
         SubCellInst_LFInst_12_LFInst_0_n9, SubCellInst_LFInst_12_LFInst_1_n26,
         SubCellInst_LFInst_12_LFInst_1_n25,
         SubCellInst_LFInst_12_LFInst_1_n24,
         SubCellInst_LFInst_12_LFInst_1_n23,
         SubCellInst_LFInst_12_LFInst_1_n22,
         SubCellInst_LFInst_12_LFInst_1_n21,
         SubCellInst_LFInst_12_LFInst_1_n20,
         SubCellInst_LFInst_12_LFInst_1_n19,
         SubCellInst_LFInst_12_LFInst_1_n18,
         SubCellInst_LFInst_12_LFInst_2_n28,
         SubCellInst_LFInst_12_LFInst_2_n27,
         SubCellInst_LFInst_12_LFInst_2_n26,
         SubCellInst_LFInst_12_LFInst_2_n25,
         SubCellInst_LFInst_12_LFInst_2_n24,
         SubCellInst_LFInst_12_LFInst_2_n23,
         SubCellInst_LFInst_12_LFInst_2_n22,
         SubCellInst_LFInst_12_LFInst_3_n26,
         SubCellInst_LFInst_12_LFInst_3_n25,
         SubCellInst_LFInst_12_LFInst_3_n24,
         SubCellInst_LFInst_12_LFInst_3_n23,
         SubCellInst_LFInst_12_LFInst_3_n22,
         SubCellInst_LFInst_12_LFInst_3_n21,
         SubCellInst_LFInst_12_LFInst_3_n20,
         SubCellInst_LFInst_12_LFInst_3_n19, SubCellInst_LFInst_13_LFInst_0_n8,
         SubCellInst_LFInst_13_LFInst_0_n7, SubCellInst_LFInst_13_LFInst_0_n6,
         SubCellInst_LFInst_13_LFInst_0_n9, SubCellInst_LFInst_13_LFInst_1_n26,
         SubCellInst_LFInst_13_LFInst_1_n25,
         SubCellInst_LFInst_13_LFInst_1_n24,
         SubCellInst_LFInst_13_LFInst_1_n23,
         SubCellInst_LFInst_13_LFInst_1_n22,
         SubCellInst_LFInst_13_LFInst_1_n21,
         SubCellInst_LFInst_13_LFInst_1_n20,
         SubCellInst_LFInst_13_LFInst_1_n19,
         SubCellInst_LFInst_13_LFInst_1_n18,
         SubCellInst_LFInst_13_LFInst_2_n29,
         SubCellInst_LFInst_13_LFInst_2_n28,
         SubCellInst_LFInst_13_LFInst_2_n27,
         SubCellInst_LFInst_13_LFInst_2_n26,
         SubCellInst_LFInst_13_LFInst_2_n25,
         SubCellInst_LFInst_13_LFInst_2_n24,
         SubCellInst_LFInst_13_LFInst_2_n23,
         SubCellInst_LFInst_13_LFInst_2_n22,
         SubCellInst_LFInst_13_LFInst_3_n26,
         SubCellInst_LFInst_13_LFInst_3_n25,
         SubCellInst_LFInst_13_LFInst_3_n24,
         SubCellInst_LFInst_13_LFInst_3_n23,
         SubCellInst_LFInst_13_LFInst_3_n22,
         SubCellInst_LFInst_13_LFInst_3_n21,
         SubCellInst_LFInst_13_LFInst_3_n20,
         SubCellInst_LFInst_13_LFInst_3_n19, SubCellInst_LFInst_14_LFInst_0_n8,
         SubCellInst_LFInst_14_LFInst_0_n7, SubCellInst_LFInst_14_LFInst_0_n6,
         SubCellInst_LFInst_14_LFInst_0_n9, SubCellInst_LFInst_14_LFInst_1_n26,
         SubCellInst_LFInst_14_LFInst_1_n25,
         SubCellInst_LFInst_14_LFInst_1_n24,
         SubCellInst_LFInst_14_LFInst_1_n23,
         SubCellInst_LFInst_14_LFInst_1_n22,
         SubCellInst_LFInst_14_LFInst_1_n21,
         SubCellInst_LFInst_14_LFInst_1_n20,
         SubCellInst_LFInst_14_LFInst_1_n19,
         SubCellInst_LFInst_14_LFInst_1_n18,
         SubCellInst_LFInst_14_LFInst_2_n28,
         SubCellInst_LFInst_14_LFInst_2_n27,
         SubCellInst_LFInst_14_LFInst_2_n26,
         SubCellInst_LFInst_14_LFInst_2_n25,
         SubCellInst_LFInst_14_LFInst_2_n24,
         SubCellInst_LFInst_14_LFInst_2_n23,
         SubCellInst_LFInst_14_LFInst_2_n22,
         SubCellInst_LFInst_14_LFInst_3_n26,
         SubCellInst_LFInst_14_LFInst_3_n25,
         SubCellInst_LFInst_14_LFInst_3_n24,
         SubCellInst_LFInst_14_LFInst_3_n23,
         SubCellInst_LFInst_14_LFInst_3_n22,
         SubCellInst_LFInst_14_LFInst_3_n21,
         SubCellInst_LFInst_14_LFInst_3_n20,
         SubCellInst_LFInst_14_LFInst_3_n19, SubCellInst_LFInst_15_LFInst_0_n8,
         SubCellInst_LFInst_15_LFInst_0_n7, SubCellInst_LFInst_15_LFInst_0_n6,
         SubCellInst_LFInst_15_LFInst_0_n9, SubCellInst_LFInst_15_LFInst_1_n26,
         SubCellInst_LFInst_15_LFInst_1_n25,
         SubCellInst_LFInst_15_LFInst_1_n24,
         SubCellInst_LFInst_15_LFInst_1_n23,
         SubCellInst_LFInst_15_LFInst_1_n22,
         SubCellInst_LFInst_15_LFInst_1_n21,
         SubCellInst_LFInst_15_LFInst_1_n20,
         SubCellInst_LFInst_15_LFInst_1_n19,
         SubCellInst_LFInst_15_LFInst_1_n18,
         SubCellInst_LFInst_15_LFInst_2_n28,
         SubCellInst_LFInst_15_LFInst_2_n27,
         SubCellInst_LFInst_15_LFInst_2_n26,
         SubCellInst_LFInst_15_LFInst_2_n25,
         SubCellInst_LFInst_15_LFInst_2_n24,
         SubCellInst_LFInst_15_LFInst_2_n23,
         SubCellInst_LFInst_15_LFInst_2_n22,
         SubCellInst_LFInst_15_LFInst_3_n26,
         SubCellInst_LFInst_15_LFInst_3_n25,
         SubCellInst_LFInst_15_LFInst_3_n24,
         SubCellInst_LFInst_15_LFInst_3_n23,
         SubCellInst_LFInst_15_LFInst_3_n22,
         SubCellInst_LFInst_15_LFInst_3_n21,
         SubCellInst_LFInst_15_LFInst_3_n20,
         SubCellInst_LFInst_15_LFInst_3_n19, MCInst_MC0_v1_0_0_,
         MCInst_MC0_v0_2Inst_0_n3, MCInst_MC0_v1_2Inst_0_n3,
         MCInst_MC0_v2_3Inst_0_n6, MCInst_MC0_v2_3Inst_0_n5,
         MCInst_MC0_v3_3Inst_0_n3, MCInst_MC0_v0_2Inst_1_n3,
         MCInst_MC0_v2_1Inst_1_n3, MCInst_MC0_v2_2Inst_1_n6,
         MCInst_MC0_v2_2Inst_1_n5, MCInst_MC0_v3_3Inst_1_n3,
         MCInst_MC0_v1_1Inst_2_n3, MCInst_MC0_v1_2Inst_2_n3,
         MCInst_MC0_v2_1Inst_2_n3, MCInst_MC0_v2_2Inst_2_n3,
         MCInst_MC0_v3_1Inst_2_n3, MCInst_MC0_v1_2Inst_3_n6,
         MCInst_MC0_v1_2Inst_3_n5, MCInst_MC0_v2_2Inst_3_n3,
         MCInst_MC0_v2_3Inst_3_n3, MCInst_MC0_r0Inst_XORInst_0_0_n8,
         MCInst_MC0_r0Inst_XORInst_0_0_n7, MCInst_MC0_r0Inst_XORInst_0_1_n8,
         MCInst_MC0_r0Inst_XORInst_0_1_n7, MCInst_MC0_r0Inst_XORInst_0_2_n8,
         MCInst_MC0_r0Inst_XORInst_0_2_n7, MCInst_MC0_r0Inst_XORInst_0_3_n8,
         MCInst_MC0_r0Inst_XORInst_0_3_n7, MCInst_MC0_r1Inst_XORInst_0_0_n8,
         MCInst_MC0_r1Inst_XORInst_0_0_n7, MCInst_MC0_r1Inst_XORInst_0_1_n8,
         MCInst_MC0_r1Inst_XORInst_0_1_n7, MCInst_MC0_r1Inst_XORInst_0_2_n8,
         MCInst_MC0_r1Inst_XORInst_0_2_n7, MCInst_MC0_r1Inst_XORInst_0_3_n8,
         MCInst_MC0_r1Inst_XORInst_0_3_n7, MCInst_MC0_r2Inst_XORInst_0_0_n8,
         MCInst_MC0_r2Inst_XORInst_0_0_n7, MCInst_MC0_r2Inst_XORInst_0_1_n8,
         MCInst_MC0_r2Inst_XORInst_0_1_n7, MCInst_MC0_r2Inst_XORInst_0_2_n8,
         MCInst_MC0_r2Inst_XORInst_0_2_n7, MCInst_MC0_r2Inst_XORInst_0_3_n8,
         MCInst_MC0_r2Inst_XORInst_0_3_n7, MCInst_MC0_r3Inst_XORInst_0_0_n8,
         MCInst_MC0_r3Inst_XORInst_0_0_n7, MCInst_MC0_r3Inst_XORInst_0_1_n8,
         MCInst_MC0_r3Inst_XORInst_0_1_n7, MCInst_MC0_r3Inst_XORInst_0_2_n8,
         MCInst_MC0_r3Inst_XORInst_0_2_n7, MCInst_MC0_r3Inst_XORInst_0_3_n8,
         MCInst_MC0_r3Inst_XORInst_0_3_n7, MCInst_MC1_v1_0_0_,
         MCInst_MC1_v0_2Inst_0_n3, MCInst_MC1_v1_2Inst_0_n3,
         MCInst_MC1_v2_3Inst_0_n6, MCInst_MC1_v2_3Inst_0_n5,
         MCInst_MC1_v3_3Inst_0_n3, MCInst_MC1_v0_2Inst_1_n3,
         MCInst_MC1_v2_1Inst_1_n3, MCInst_MC1_v2_2Inst_1_n6,
         MCInst_MC1_v2_2Inst_1_n5, MCInst_MC1_v3_3Inst_1_n3,
         MCInst_MC1_v1_1Inst_2_n3, MCInst_MC1_v1_2Inst_2_n3,
         MCInst_MC1_v2_1Inst_2_n3, MCInst_MC1_v2_2Inst_2_n3,
         MCInst_MC1_v3_1Inst_2_n3, MCInst_MC1_v1_2Inst_3_n6,
         MCInst_MC1_v1_2Inst_3_n5, MCInst_MC1_v2_2Inst_3_n3,
         MCInst_MC1_v2_3Inst_3_n3, MCInst_MC1_r0Inst_XORInst_0_0_n8,
         MCInst_MC1_r0Inst_XORInst_0_0_n7, MCInst_MC1_r0Inst_XORInst_0_1_n8,
         MCInst_MC1_r0Inst_XORInst_0_1_n7, MCInst_MC1_r0Inst_XORInst_0_2_n8,
         MCInst_MC1_r0Inst_XORInst_0_2_n7, MCInst_MC1_r0Inst_XORInst_0_3_n8,
         MCInst_MC1_r0Inst_XORInst_0_3_n7, MCInst_MC1_r1Inst_XORInst_0_0_n8,
         MCInst_MC1_r1Inst_XORInst_0_0_n7, MCInst_MC1_r1Inst_XORInst_0_1_n8,
         MCInst_MC1_r1Inst_XORInst_0_1_n7, MCInst_MC1_r1Inst_XORInst_0_2_n8,
         MCInst_MC1_r1Inst_XORInst_0_2_n7, MCInst_MC1_r1Inst_XORInst_0_3_n8,
         MCInst_MC1_r1Inst_XORInst_0_3_n7, MCInst_MC1_r2Inst_XORInst_0_0_n8,
         MCInst_MC1_r2Inst_XORInst_0_0_n7, MCInst_MC1_r2Inst_XORInst_0_1_n8,
         MCInst_MC1_r2Inst_XORInst_0_1_n7, MCInst_MC1_r2Inst_XORInst_0_2_n8,
         MCInst_MC1_r2Inst_XORInst_0_2_n7, MCInst_MC1_r2Inst_XORInst_0_3_n8,
         MCInst_MC1_r2Inst_XORInst_0_3_n7, MCInst_MC1_r3Inst_XORInst_0_0_n8,
         MCInst_MC1_r3Inst_XORInst_0_0_n7, MCInst_MC1_r3Inst_XORInst_0_1_n8,
         MCInst_MC1_r3Inst_XORInst_0_1_n7, MCInst_MC1_r3Inst_XORInst_0_2_n8,
         MCInst_MC1_r3Inst_XORInst_0_2_n7, MCInst_MC1_r3Inst_XORInst_0_3_n8,
         MCInst_MC1_r3Inst_XORInst_0_3_n7, MCInst_MC2_v1_0_0_,
         MCInst_MC2_v0_2Inst_0_n3, MCInst_MC2_v1_2Inst_0_n3,
         MCInst_MC2_v2_3Inst_0_n6, MCInst_MC2_v2_3Inst_0_n5,
         MCInst_MC2_v3_3Inst_0_n3, MCInst_MC2_v0_2Inst_1_n3,
         MCInst_MC2_v2_1Inst_1_n3, MCInst_MC2_v2_2Inst_1_n6,
         MCInst_MC2_v2_2Inst_1_n5, MCInst_MC2_v3_3Inst_1_n3,
         MCInst_MC2_v1_1Inst_2_n3, MCInst_MC2_v1_2Inst_2_n3,
         MCInst_MC2_v2_1Inst_2_n3, MCInst_MC2_v2_2Inst_2_n3,
         MCInst_MC2_v3_1Inst_2_n3, MCInst_MC2_v1_2Inst_3_n6,
         MCInst_MC2_v1_2Inst_3_n5, MCInst_MC2_v2_2Inst_3_n3,
         MCInst_MC2_v2_3Inst_3_n3, MCInst_MC2_r0Inst_XORInst_0_0_n8,
         MCInst_MC2_r0Inst_XORInst_0_0_n7, MCInst_MC2_r0Inst_XORInst_0_1_n8,
         MCInst_MC2_r0Inst_XORInst_0_1_n7, MCInst_MC2_r0Inst_XORInst_0_2_n8,
         MCInst_MC2_r0Inst_XORInst_0_2_n7, MCInst_MC2_r0Inst_XORInst_0_3_n8,
         MCInst_MC2_r0Inst_XORInst_0_3_n7, MCInst_MC2_r1Inst_XORInst_0_0_n8,
         MCInst_MC2_r1Inst_XORInst_0_0_n7, MCInst_MC2_r1Inst_XORInst_0_1_n8,
         MCInst_MC2_r1Inst_XORInst_0_1_n7, MCInst_MC2_r1Inst_XORInst_0_2_n8,
         MCInst_MC2_r1Inst_XORInst_0_2_n7, MCInst_MC2_r1Inst_XORInst_0_3_n8,
         MCInst_MC2_r1Inst_XORInst_0_3_n7, MCInst_MC2_r2Inst_XORInst_0_0_n8,
         MCInst_MC2_r2Inst_XORInst_0_0_n7, MCInst_MC2_r2Inst_XORInst_0_1_n8,
         MCInst_MC2_r2Inst_XORInst_0_1_n7, MCInst_MC2_r2Inst_XORInst_0_2_n8,
         MCInst_MC2_r2Inst_XORInst_0_2_n7, MCInst_MC2_r2Inst_XORInst_0_3_n8,
         MCInst_MC2_r2Inst_XORInst_0_3_n7, MCInst_MC2_r3Inst_XORInst_0_0_n8,
         MCInst_MC2_r3Inst_XORInst_0_0_n7, MCInst_MC2_r3Inst_XORInst_0_1_n8,
         MCInst_MC2_r3Inst_XORInst_0_1_n7, MCInst_MC2_r3Inst_XORInst_0_2_n8,
         MCInst_MC2_r3Inst_XORInst_0_2_n7, MCInst_MC2_r3Inst_XORInst_0_3_n8,
         MCInst_MC2_r3Inst_XORInst_0_3_n7, MCInst_MC3_v1_0_0_,
         MCInst_MC3_v0_2Inst_0_n3, MCInst_MC3_v1_2Inst_0_n3,
         MCInst_MC3_v2_3Inst_0_n6, MCInst_MC3_v2_3Inst_0_n5,
         MCInst_MC3_v3_3Inst_0_n3, MCInst_MC3_v0_2Inst_1_n3,
         MCInst_MC3_v2_1Inst_1_n3, MCInst_MC3_v2_2Inst_1_n6,
         MCInst_MC3_v2_2Inst_1_n5, MCInst_MC3_v3_3Inst_1_n3,
         MCInst_MC3_v1_1Inst_2_n3, MCInst_MC3_v1_2Inst_2_n3,
         MCInst_MC3_v2_1Inst_2_n3, MCInst_MC3_v2_2Inst_2_n3,
         MCInst_MC3_v3_1Inst_2_n3, MCInst_MC3_v1_2Inst_3_n6,
         MCInst_MC3_v1_2Inst_3_n5, MCInst_MC3_v2_2Inst_3_n3,
         MCInst_MC3_v2_3Inst_3_n3, MCInst_MC3_r0Inst_XORInst_0_0_n8,
         MCInst_MC3_r0Inst_XORInst_0_0_n7, MCInst_MC3_r0Inst_XORInst_0_1_n8,
         MCInst_MC3_r0Inst_XORInst_0_1_n7, MCInst_MC3_r0Inst_XORInst_0_2_n8,
         MCInst_MC3_r0Inst_XORInst_0_2_n7, MCInst_MC3_r0Inst_XORInst_0_3_n8,
         MCInst_MC3_r0Inst_XORInst_0_3_n7, MCInst_MC3_r1Inst_XORInst_0_0_n8,
         MCInst_MC3_r1Inst_XORInst_0_0_n7, MCInst_MC3_r1Inst_XORInst_0_1_n8,
         MCInst_MC3_r1Inst_XORInst_0_1_n7, MCInst_MC3_r1Inst_XORInst_0_2_n8,
         MCInst_MC3_r1Inst_XORInst_0_2_n7, MCInst_MC3_r1Inst_XORInst_0_3_n8,
         MCInst_MC3_r1Inst_XORInst_0_3_n7, MCInst_MC3_r2Inst_XORInst_0_0_n8,
         MCInst_MC3_r2Inst_XORInst_0_0_n7, MCInst_MC3_r2Inst_XORInst_0_1_n8,
         MCInst_MC3_r2Inst_XORInst_0_1_n7, MCInst_MC3_r2Inst_XORInst_0_2_n8,
         MCInst_MC3_r2Inst_XORInst_0_2_n7, MCInst_MC3_r2Inst_XORInst_0_3_n8,
         MCInst_MC3_r2Inst_XORInst_0_3_n7, MCInst_MC3_r3Inst_XORInst_0_0_n8,
         MCInst_MC3_r3Inst_XORInst_0_0_n7, MCInst_MC3_r3Inst_XORInst_0_1_n8,
         MCInst_MC3_r3Inst_XORInst_0_1_n7, MCInst_MC3_r3Inst_XORInst_0_2_n8,
         MCInst_MC3_r3Inst_XORInst_0_2_n7, MCInst_MC3_r3Inst_XORInst_0_3_n8,
         MCInst_MC3_r3Inst_XORInst_0_3_n7,
         Red_PlaintextInst_LFInst_0_LFInst_0_n3,
         Red_PlaintextInst_LFInst_0_LFInst_1_n3,
         Red_PlaintextInst_LFInst_0_LFInst_2_n3,
         Red_PlaintextInst_LFInst_1_LFInst_0_n3,
         Red_PlaintextInst_LFInst_1_LFInst_1_n3,
         Red_PlaintextInst_LFInst_1_LFInst_2_n3,
         Red_PlaintextInst_LFInst_2_LFInst_0_n3,
         Red_PlaintextInst_LFInst_2_LFInst_1_n3,
         Red_PlaintextInst_LFInst_2_LFInst_2_n3,
         Red_PlaintextInst_LFInst_3_LFInst_0_n3,
         Red_PlaintextInst_LFInst_3_LFInst_1_n3,
         Red_PlaintextInst_LFInst_3_LFInst_2_n3,
         Red_PlaintextInst_LFInst_4_LFInst_0_n3,
         Red_PlaintextInst_LFInst_4_LFInst_1_n3,
         Red_PlaintextInst_LFInst_4_LFInst_2_n3,
         Red_PlaintextInst_LFInst_5_LFInst_0_n3,
         Red_PlaintextInst_LFInst_5_LFInst_1_n3,
         Red_PlaintextInst_LFInst_5_LFInst_2_n3,
         Red_PlaintextInst_LFInst_6_LFInst_0_n3,
         Red_PlaintextInst_LFInst_6_LFInst_1_n3,
         Red_PlaintextInst_LFInst_6_LFInst_2_n3,
         Red_PlaintextInst_LFInst_7_LFInst_0_n3,
         Red_PlaintextInst_LFInst_7_LFInst_1_n3,
         Red_PlaintextInst_LFInst_7_LFInst_2_n3,
         Red_PlaintextInst_LFInst_8_LFInst_0_n3,
         Red_PlaintextInst_LFInst_8_LFInst_1_n3,
         Red_PlaintextInst_LFInst_8_LFInst_2_n3,
         Red_PlaintextInst_LFInst_9_LFInst_0_n3,
         Red_PlaintextInst_LFInst_9_LFInst_1_n3,
         Red_PlaintextInst_LFInst_9_LFInst_2_n3,
         Red_PlaintextInst_LFInst_10_LFInst_0_n3,
         Red_PlaintextInst_LFInst_10_LFInst_1_n3,
         Red_PlaintextInst_LFInst_10_LFInst_2_n3,
         Red_PlaintextInst_LFInst_11_LFInst_0_n3,
         Red_PlaintextInst_LFInst_11_LFInst_1_n3,
         Red_PlaintextInst_LFInst_11_LFInst_2_n3,
         Red_PlaintextInst_LFInst_12_LFInst_0_n3,
         Red_PlaintextInst_LFInst_12_LFInst_1_n3,
         Red_PlaintextInst_LFInst_12_LFInst_2_n3,
         Red_PlaintextInst_LFInst_13_LFInst_0_n3,
         Red_PlaintextInst_LFInst_13_LFInst_1_n3,
         Red_PlaintextInst_LFInst_13_LFInst_2_n3,
         Red_PlaintextInst_LFInst_14_LFInst_0_n3,
         Red_PlaintextInst_LFInst_14_LFInst_1_n3,
         Red_PlaintextInst_LFInst_14_LFInst_2_n3,
         Red_PlaintextInst_LFInst_15_LFInst_0_n3,
         Red_PlaintextInst_LFInst_15_LFInst_1_n3,
         Red_PlaintextInst_LFInst_15_LFInst_2_n3,
         Red_SubCellInst_LFInst_0_LFInst_0_n12,
         Red_SubCellInst_LFInst_0_LFInst_0_n11,
         Red_SubCellInst_LFInst_0_LFInst_0_n10,
         Red_SubCellInst_LFInst_0_LFInst_0_n9,
         Red_SubCellInst_LFInst_0_LFInst_1_n6,
         Red_SubCellInst_LFInst_0_LFInst_1_n5,
         Red_SubCellInst_LFInst_0_LFInst_2_n17,
         Red_SubCellInst_LFInst_0_LFInst_2_n16,
         Red_SubCellInst_LFInst_0_LFInst_2_n15,
         Red_SubCellInst_LFInst_0_LFInst_2_n14,
         Red_SubCellInst_LFInst_0_LFInst_2_n13,
         Red_SubCellInst_LFInst_0_LFInst_2_n12,
         Red_SubCellInst_LFInst_1_LFInst_0_n12,
         Red_SubCellInst_LFInst_1_LFInst_0_n11,
         Red_SubCellInst_LFInst_1_LFInst_0_n10,
         Red_SubCellInst_LFInst_1_LFInst_0_n9,
         Red_SubCellInst_LFInst_1_LFInst_1_n6,
         Red_SubCellInst_LFInst_1_LFInst_1_n5,
         Red_SubCellInst_LFInst_1_LFInst_2_n16,
         Red_SubCellInst_LFInst_1_LFInst_2_n15,
         Red_SubCellInst_LFInst_1_LFInst_2_n14,
         Red_SubCellInst_LFInst_1_LFInst_2_n13,
         Red_SubCellInst_LFInst_1_LFInst_2_n12,
         Red_SubCellInst_LFInst_2_LFInst_0_n12,
         Red_SubCellInst_LFInst_2_LFInst_0_n11,
         Red_SubCellInst_LFInst_2_LFInst_0_n10,
         Red_SubCellInst_LFInst_2_LFInst_0_n9,
         Red_SubCellInst_LFInst_2_LFInst_1_n6,
         Red_SubCellInst_LFInst_2_LFInst_1_n5,
         Red_SubCellInst_LFInst_2_LFInst_2_n16,
         Red_SubCellInst_LFInst_2_LFInst_2_n15,
         Red_SubCellInst_LFInst_2_LFInst_2_n14,
         Red_SubCellInst_LFInst_2_LFInst_2_n13,
         Red_SubCellInst_LFInst_2_LFInst_2_n12,
         Red_SubCellInst_LFInst_3_LFInst_0_n12,
         Red_SubCellInst_LFInst_3_LFInst_0_n11,
         Red_SubCellInst_LFInst_3_LFInst_0_n10,
         Red_SubCellInst_LFInst_3_LFInst_0_n9,
         Red_SubCellInst_LFInst_3_LFInst_1_n6,
         Red_SubCellInst_LFInst_3_LFInst_1_n5,
         Red_SubCellInst_LFInst_3_LFInst_2_n16,
         Red_SubCellInst_LFInst_3_LFInst_2_n15,
         Red_SubCellInst_LFInst_3_LFInst_2_n14,
         Red_SubCellInst_LFInst_3_LFInst_2_n13,
         Red_SubCellInst_LFInst_3_LFInst_2_n12,
         Red_SubCellInst_LFInst_4_LFInst_0_n12,
         Red_SubCellInst_LFInst_4_LFInst_0_n11,
         Red_SubCellInst_LFInst_4_LFInst_0_n10,
         Red_SubCellInst_LFInst_4_LFInst_0_n9,
         Red_SubCellInst_LFInst_4_LFInst_1_n6,
         Red_SubCellInst_LFInst_4_LFInst_1_n5,
         Red_SubCellInst_LFInst_4_LFInst_2_n16,
         Red_SubCellInst_LFInst_4_LFInst_2_n15,
         Red_SubCellInst_LFInst_4_LFInst_2_n14,
         Red_SubCellInst_LFInst_4_LFInst_2_n13,
         Red_SubCellInst_LFInst_4_LFInst_2_n12,
         Red_SubCellInst_LFInst_5_LFInst_0_n12,
         Red_SubCellInst_LFInst_5_LFInst_0_n11,
         Red_SubCellInst_LFInst_5_LFInst_0_n10,
         Red_SubCellInst_LFInst_5_LFInst_0_n9,
         Red_SubCellInst_LFInst_5_LFInst_1_n6,
         Red_SubCellInst_LFInst_5_LFInst_1_n5,
         Red_SubCellInst_LFInst_5_LFInst_2_n16,
         Red_SubCellInst_LFInst_5_LFInst_2_n15,
         Red_SubCellInst_LFInst_5_LFInst_2_n14,
         Red_SubCellInst_LFInst_5_LFInst_2_n13,
         Red_SubCellInst_LFInst_5_LFInst_2_n12,
         Red_SubCellInst_LFInst_6_LFInst_0_n12,
         Red_SubCellInst_LFInst_6_LFInst_0_n11,
         Red_SubCellInst_LFInst_6_LFInst_0_n10,
         Red_SubCellInst_LFInst_6_LFInst_0_n9,
         Red_SubCellInst_LFInst_6_LFInst_1_n6,
         Red_SubCellInst_LFInst_6_LFInst_1_n5,
         Red_SubCellInst_LFInst_6_LFInst_2_n16,
         Red_SubCellInst_LFInst_6_LFInst_2_n15,
         Red_SubCellInst_LFInst_6_LFInst_2_n14,
         Red_SubCellInst_LFInst_6_LFInst_2_n13,
         Red_SubCellInst_LFInst_6_LFInst_2_n12,
         Red_SubCellInst_LFInst_7_LFInst_0_n12,
         Red_SubCellInst_LFInst_7_LFInst_0_n11,
         Red_SubCellInst_LFInst_7_LFInst_0_n10,
         Red_SubCellInst_LFInst_7_LFInst_0_n9,
         Red_SubCellInst_LFInst_7_LFInst_1_n6,
         Red_SubCellInst_LFInst_7_LFInst_1_n5,
         Red_SubCellInst_LFInst_7_LFInst_2_n17,
         Red_SubCellInst_LFInst_7_LFInst_2_n16,
         Red_SubCellInst_LFInst_7_LFInst_2_n15,
         Red_SubCellInst_LFInst_7_LFInst_2_n14,
         Red_SubCellInst_LFInst_7_LFInst_2_n13,
         Red_SubCellInst_LFInst_7_LFInst_2_n12,
         Red_SubCellInst_LFInst_8_LFInst_0_n12,
         Red_SubCellInst_LFInst_8_LFInst_0_n11,
         Red_SubCellInst_LFInst_8_LFInst_0_n10,
         Red_SubCellInst_LFInst_8_LFInst_0_n9,
         Red_SubCellInst_LFInst_8_LFInst_1_n6,
         Red_SubCellInst_LFInst_8_LFInst_1_n5,
         Red_SubCellInst_LFInst_8_LFInst_2_n16,
         Red_SubCellInst_LFInst_8_LFInst_2_n15,
         Red_SubCellInst_LFInst_8_LFInst_2_n14,
         Red_SubCellInst_LFInst_8_LFInst_2_n13,
         Red_SubCellInst_LFInst_8_LFInst_2_n12,
         Red_SubCellInst_LFInst_9_LFInst_0_n12,
         Red_SubCellInst_LFInst_9_LFInst_0_n11,
         Red_SubCellInst_LFInst_9_LFInst_0_n10,
         Red_SubCellInst_LFInst_9_LFInst_0_n9,
         Red_SubCellInst_LFInst_9_LFInst_1_n6,
         Red_SubCellInst_LFInst_9_LFInst_1_n5,
         Red_SubCellInst_LFInst_9_LFInst_2_n13,
         Red_SubCellInst_LFInst_9_LFInst_2_n12,
         Red_SubCellInst_LFInst_9_LFInst_2_n11,
         Red_SubCellInst_LFInst_9_LFInst_2_n10,
         Red_SubCellInst_LFInst_9_LFInst_2_n9,
         Red_SubCellInst_LFInst_10_LFInst_0_n12,
         Red_SubCellInst_LFInst_10_LFInst_0_n11,
         Red_SubCellInst_LFInst_10_LFInst_0_n10,
         Red_SubCellInst_LFInst_10_LFInst_0_n9,
         Red_SubCellInst_LFInst_10_LFInst_1_n6,
         Red_SubCellInst_LFInst_10_LFInst_1_n5,
         Red_SubCellInst_LFInst_10_LFInst_2_n16,
         Red_SubCellInst_LFInst_10_LFInst_2_n15,
         Red_SubCellInst_LFInst_10_LFInst_2_n14,
         Red_SubCellInst_LFInst_10_LFInst_2_n13,
         Red_SubCellInst_LFInst_10_LFInst_2_n12,
         Red_SubCellInst_LFInst_11_LFInst_0_n12,
         Red_SubCellInst_LFInst_11_LFInst_0_n11,
         Red_SubCellInst_LFInst_11_LFInst_0_n10,
         Red_SubCellInst_LFInst_11_LFInst_0_n9,
         Red_SubCellInst_LFInst_11_LFInst_1_n6,
         Red_SubCellInst_LFInst_11_LFInst_1_n5,
         Red_SubCellInst_LFInst_11_LFInst_2_n17,
         Red_SubCellInst_LFInst_11_LFInst_2_n16,
         Red_SubCellInst_LFInst_11_LFInst_2_n15,
         Red_SubCellInst_LFInst_11_LFInst_2_n14,
         Red_SubCellInst_LFInst_11_LFInst_2_n13,
         Red_SubCellInst_LFInst_11_LFInst_2_n12,
         Red_SubCellInst_LFInst_12_LFInst_0_n12,
         Red_SubCellInst_LFInst_12_LFInst_0_n11,
         Red_SubCellInst_LFInst_12_LFInst_0_n10,
         Red_SubCellInst_LFInst_12_LFInst_0_n9,
         Red_SubCellInst_LFInst_12_LFInst_1_n6,
         Red_SubCellInst_LFInst_12_LFInst_1_n5,
         Red_SubCellInst_LFInst_12_LFInst_2_n16,
         Red_SubCellInst_LFInst_12_LFInst_2_n15,
         Red_SubCellInst_LFInst_12_LFInst_2_n14,
         Red_SubCellInst_LFInst_12_LFInst_2_n13,
         Red_SubCellInst_LFInst_12_LFInst_2_n12,
         Red_SubCellInst_LFInst_13_LFInst_0_n12,
         Red_SubCellInst_LFInst_13_LFInst_0_n11,
         Red_SubCellInst_LFInst_13_LFInst_0_n10,
         Red_SubCellInst_LFInst_13_LFInst_0_n9,
         Red_SubCellInst_LFInst_13_LFInst_1_n6,
         Red_SubCellInst_LFInst_13_LFInst_1_n5,
         Red_SubCellInst_LFInst_13_LFInst_2_n16,
         Red_SubCellInst_LFInst_13_LFInst_2_n15,
         Red_SubCellInst_LFInst_13_LFInst_2_n14,
         Red_SubCellInst_LFInst_13_LFInst_2_n13,
         Red_SubCellInst_LFInst_13_LFInst_2_n12,
         Red_SubCellInst_LFInst_14_LFInst_0_n12,
         Red_SubCellInst_LFInst_14_LFInst_0_n11,
         Red_SubCellInst_LFInst_14_LFInst_0_n10,
         Red_SubCellInst_LFInst_14_LFInst_0_n9,
         Red_SubCellInst_LFInst_14_LFInst_1_n6,
         Red_SubCellInst_LFInst_14_LFInst_1_n5,
         Red_SubCellInst_LFInst_14_LFInst_2_n16,
         Red_SubCellInst_LFInst_14_LFInst_2_n15,
         Red_SubCellInst_LFInst_14_LFInst_2_n14,
         Red_SubCellInst_LFInst_14_LFInst_2_n13,
         Red_SubCellInst_LFInst_14_LFInst_2_n12,
         Red_SubCellInst_LFInst_15_LFInst_0_n12,
         Red_SubCellInst_LFInst_15_LFInst_0_n11,
         Red_SubCellInst_LFInst_15_LFInst_0_n10,
         Red_SubCellInst_LFInst_15_LFInst_0_n9,
         Red_SubCellInst_LFInst_15_LFInst_1_n6,
         Red_SubCellInst_LFInst_15_LFInst_1_n5,
         Red_SubCellInst_LFInst_15_LFInst_2_n16,
         Red_SubCellInst_LFInst_15_LFInst_2_n15,
         Red_SubCellInst_LFInst_15_LFInst_2_n14,
         Red_SubCellInst_LFInst_15_LFInst_2_n13,
         Red_SubCellInst_LFInst_15_LFInst_2_n12, Red_MCInst_MC0_v1_0Inst_0_n3,
         Red_MCInst_MC0_v2_2Inst_0_n3, Red_MCInst_MC0_v2_3Inst_0_n3,
         Red_MCInst_MC0_v3_2Inst_0_n6, Red_MCInst_MC0_v3_2Inst_0_n5,
         Red_MCInst_MC0_v0_1Inst_1_n3, Red_MCInst_MC0_v1_0Inst_1_n3,
         Red_MCInst_MC0_v1_1Inst_1_n6, Red_MCInst_MC0_v1_1Inst_1_n5,
         Red_MCInst_MC0_v3_1Inst_1_n6, Red_MCInst_MC0_v3_1Inst_1_n5,
         Red_MCInst_MC0_v0_0Inst_2_n3, Red_MCInst_MC0_v0_3Inst_2_n6,
         Red_MCInst_MC0_v0_3Inst_2_n5, Red_MCInst_MC0_v1_0Inst_2_n3,
         Red_MCInst_MC0_v1_2Inst_2_n3, Red_MCInst_MC0_v1_3Inst_2_n6,
         Red_MCInst_MC0_v1_3Inst_2_n5, Red_MCInst_MC0_v2_0Inst_2_n6,
         Red_MCInst_MC0_v2_0Inst_2_n5, Red_MCInst_MC0_v3_0Inst_2_n6,
         Red_MCInst_MC0_v3_0Inst_2_n5, Red_MCInst_MC0_v3_2Inst_2_n3,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_2_n7, Red_MCInst_MC1_v1_0Inst_0_n3,
         Red_MCInst_MC1_v2_2Inst_0_n3, Red_MCInst_MC1_v2_3Inst_0_n3,
         Red_MCInst_MC1_v3_2Inst_0_n6, Red_MCInst_MC1_v3_2Inst_0_n5,
         Red_MCInst_MC1_v0_1Inst_1_n3, Red_MCInst_MC1_v1_0Inst_1_n3,
         Red_MCInst_MC1_v1_1Inst_1_n6, Red_MCInst_MC1_v1_1Inst_1_n5,
         Red_MCInst_MC1_v3_1Inst_1_n6, Red_MCInst_MC1_v3_1Inst_1_n5,
         Red_MCInst_MC1_v0_0Inst_2_n3, Red_MCInst_MC1_v0_3Inst_2_n6,
         Red_MCInst_MC1_v0_3Inst_2_n5, Red_MCInst_MC1_v1_0Inst_2_n3,
         Red_MCInst_MC1_v1_2Inst_2_n3, Red_MCInst_MC1_v1_3Inst_2_n6,
         Red_MCInst_MC1_v1_3Inst_2_n5, Red_MCInst_MC1_v2_0Inst_2_n6,
         Red_MCInst_MC1_v2_0Inst_2_n5, Red_MCInst_MC1_v3_0Inst_2_n6,
         Red_MCInst_MC1_v3_0Inst_2_n5, Red_MCInst_MC1_v3_2Inst_2_n3,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_2_n7, Red_MCInst_MC2_v1_0Inst_0_n3,
         Red_MCInst_MC2_v2_2Inst_0_n3, Red_MCInst_MC2_v2_3Inst_0_n3,
         Red_MCInst_MC2_v3_2Inst_0_n6, Red_MCInst_MC2_v3_2Inst_0_n5,
         Red_MCInst_MC2_v0_1Inst_1_n3, Red_MCInst_MC2_v1_0Inst_1_n3,
         Red_MCInst_MC2_v1_1Inst_1_n6, Red_MCInst_MC2_v1_1Inst_1_n5,
         Red_MCInst_MC2_v3_1Inst_1_n6, Red_MCInst_MC2_v3_1Inst_1_n5,
         Red_MCInst_MC2_v0_0Inst_2_n3, Red_MCInst_MC2_v0_3Inst_2_n6,
         Red_MCInst_MC2_v0_3Inst_2_n5, Red_MCInst_MC2_v1_0Inst_2_n3,
         Red_MCInst_MC2_v1_2Inst_2_n3, Red_MCInst_MC2_v1_3Inst_2_n6,
         Red_MCInst_MC2_v1_3Inst_2_n5, Red_MCInst_MC2_v2_0Inst_2_n6,
         Red_MCInst_MC2_v2_0Inst_2_n5, Red_MCInst_MC2_v3_0Inst_2_n6,
         Red_MCInst_MC2_v3_0Inst_2_n5, Red_MCInst_MC2_v3_2Inst_2_n3,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_2_n7, Red_MCInst_MC3_v1_0Inst_0_n3,
         Red_MCInst_MC3_v2_2Inst_0_n3, Red_MCInst_MC3_v2_3Inst_0_n3,
         Red_MCInst_MC3_v3_2Inst_0_n6, Red_MCInst_MC3_v3_2Inst_0_n5,
         Red_MCInst_MC3_v0_1Inst_1_n3, Red_MCInst_MC3_v1_0Inst_1_n3,
         Red_MCInst_MC3_v1_1Inst_1_n6, Red_MCInst_MC3_v1_1Inst_1_n5,
         Red_MCInst_MC3_v3_1Inst_1_n6, Red_MCInst_MC3_v3_1Inst_1_n5,
         Red_MCInst_MC3_v0_0Inst_2_n3, Red_MCInst_MC3_v0_3Inst_2_n6,
         Red_MCInst_MC3_v0_3Inst_2_n5, Red_MCInst_MC3_v1_0Inst_2_n3,
         Red_MCInst_MC3_v1_2Inst_2_n3, Red_MCInst_MC3_v1_3Inst_2_n6,
         Red_MCInst_MC3_v1_3Inst_2_n5, Red_MCInst_MC3_v2_0Inst_2_n6,
         Red_MCInst_MC3_v2_0Inst_2_n5, Red_MCInst_MC3_v3_0Inst_2_n6,
         Red_MCInst_MC3_v3_0Inst_2_n5, Red_MCInst_MC3_v3_2Inst_2_n3,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_2_n7,
         Red_KeyInst_LFInst_0_LFInst_0_n3, Red_KeyInst_LFInst_0_LFInst_1_n3,
         Red_KeyInst_LFInst_0_LFInst_2_n3, Red_KeyInst_LFInst_1_LFInst_0_n3,
         Red_KeyInst_LFInst_1_LFInst_1_n3, Red_KeyInst_LFInst_1_LFInst_2_n3,
         Red_KeyInst_LFInst_2_LFInst_0_n3, Red_KeyInst_LFInst_2_LFInst_1_n3,
         Red_KeyInst_LFInst_2_LFInst_2_n3, Red_KeyInst_LFInst_3_LFInst_0_n3,
         Red_KeyInst_LFInst_3_LFInst_1_n3, Red_KeyInst_LFInst_3_LFInst_2_n3,
         Red_KeyInst_LFInst_4_LFInst_0_n3, Red_KeyInst_LFInst_4_LFInst_1_n3,
         Red_KeyInst_LFInst_4_LFInst_2_n3, Red_KeyInst_LFInst_5_LFInst_0_n3,
         Red_KeyInst_LFInst_5_LFInst_1_n3, Red_KeyInst_LFInst_5_LFInst_2_n3,
         Red_KeyInst_LFInst_6_LFInst_0_n3, Red_KeyInst_LFInst_6_LFInst_1_n3,
         Red_KeyInst_LFInst_6_LFInst_2_n3, Red_KeyInst_LFInst_7_LFInst_0_n3,
         Red_KeyInst_LFInst_7_LFInst_1_n3, Red_KeyInst_LFInst_7_LFInst_2_n3,
         Red_KeyInst_LFInst_8_LFInst_0_n3, Red_KeyInst_LFInst_8_LFInst_1_n3,
         Red_KeyInst_LFInst_8_LFInst_2_n3, Red_KeyInst_LFInst_9_LFInst_0_n3,
         Red_KeyInst_LFInst_9_LFInst_1_n3, Red_KeyInst_LFInst_9_LFInst_2_n3,
         Red_KeyInst_LFInst_10_LFInst_0_n3, Red_KeyInst_LFInst_10_LFInst_1_n3,
         Red_KeyInst_LFInst_10_LFInst_2_n3, Red_KeyInst_LFInst_11_LFInst_0_n3,
         Red_KeyInst_LFInst_11_LFInst_1_n3, Red_KeyInst_LFInst_11_LFInst_2_n3,
         Red_KeyInst_LFInst_12_LFInst_0_n3, Red_KeyInst_LFInst_12_LFInst_1_n3,
         Red_KeyInst_LFInst_12_LFInst_2_n3, Red_KeyInst_LFInst_13_LFInst_0_n3,
         Red_KeyInst_LFInst_13_LFInst_1_n3, Red_KeyInst_LFInst_13_LFInst_2_n3,
         Red_KeyInst_LFInst_14_LFInst_0_n3, Red_KeyInst_LFInst_14_LFInst_1_n3,
         Red_KeyInst_LFInst_14_LFInst_2_n3, Red_KeyInst_LFInst_15_LFInst_0_n3,
         Red_KeyInst_LFInst_15_LFInst_1_n3, Red_KeyInst_LFInst_15_LFInst_2_n3,
         Red_ToCheckInst_LFInst_0_LFInst_0_n3,
         Red_ToCheckInst_LFInst_0_LFInst_1_n3,
         Red_ToCheckInst_LFInst_0_LFInst_2_n3,
         Red_ToCheckInst_LFInst_1_LFInst_0_n3,
         Red_ToCheckInst_LFInst_1_LFInst_1_n3,
         Red_ToCheckInst_LFInst_1_LFInst_2_n3,
         Red_ToCheckInst_LFInst_2_LFInst_0_n3,
         Red_ToCheckInst_LFInst_2_LFInst_1_n3,
         Red_ToCheckInst_LFInst_2_LFInst_2_n3,
         Red_ToCheckInst_LFInst_3_LFInst_0_n3,
         Red_ToCheckInst_LFInst_3_LFInst_1_n3,
         Red_ToCheckInst_LFInst_3_LFInst_2_n3,
         Red_ToCheckInst_LFInst_4_LFInst_0_n3,
         Red_ToCheckInst_LFInst_4_LFInst_1_n3,
         Red_ToCheckInst_LFInst_4_LFInst_2_n3,
         Red_ToCheckInst_LFInst_5_LFInst_0_n3,
         Red_ToCheckInst_LFInst_5_LFInst_1_n3,
         Red_ToCheckInst_LFInst_5_LFInst_2_n3,
         Red_ToCheckInst_LFInst_6_LFInst_0_n3,
         Red_ToCheckInst_LFInst_6_LFInst_1_n3,
         Red_ToCheckInst_LFInst_6_LFInst_2_n3,
         Red_ToCheckInst_LFInst_7_LFInst_0_n3,
         Red_ToCheckInst_LFInst_7_LFInst_1_n3,
         Red_ToCheckInst_LFInst_7_LFInst_2_n3,
         Red_ToCheckInst_LFInst_8_LFInst_0_n3,
         Red_ToCheckInst_LFInst_8_LFInst_1_n3,
         Red_ToCheckInst_LFInst_8_LFInst_2_n3,
         Red_ToCheckInst_LFInst_9_LFInst_0_n3,
         Red_ToCheckInst_LFInst_9_LFInst_1_n3,
         Red_ToCheckInst_LFInst_9_LFInst_2_n3,
         Red_ToCheckInst_LFInst_10_LFInst_0_n3,
         Red_ToCheckInst_LFInst_10_LFInst_1_n3,
         Red_ToCheckInst_LFInst_10_LFInst_2_n3,
         Red_ToCheckInst_LFInst_11_LFInst_0_n3,
         Red_ToCheckInst_LFInst_11_LFInst_1_n3,
         Red_ToCheckInst_LFInst_11_LFInst_2_n3,
         Red_ToCheckInst_LFInst_12_LFInst_0_n3,
         Red_ToCheckInst_LFInst_12_LFInst_1_n3,
         Red_ToCheckInst_LFInst_12_LFInst_2_n3,
         Red_ToCheckInst_LFInst_13_LFInst_0_n3,
         Red_ToCheckInst_LFInst_13_LFInst_1_n3,
         Red_ToCheckInst_LFInst_13_LFInst_2_n3,
         Red_ToCheckInst_LFInst_14_LFInst_0_n3,
         Red_ToCheckInst_LFInst_14_LFInst_1_n3,
         Red_ToCheckInst_LFInst_14_LFInst_2_n3,
         Red_ToCheckInst_LFInst_15_LFInst_0_n3,
         Red_ToCheckInst_LFInst_15_LFInst_1_n3,
         Red_ToCheckInst_LFInst_15_LFInst_2_n3,
         Red_ToCheckInst_LFInst_16_LFInst_0_n3,
         Red_ToCheckInst_LFInst_16_LFInst_1_n3,
         Red_ToCheckInst_LFInst_16_LFInst_2_n3,
         Red_ToCheckInst_LFInst_17_LFInst_0_n3,
         Red_ToCheckInst_LFInst_17_LFInst_1_n3,
         Red_ToCheckInst_LFInst_17_LFInst_2_n3,
         Red_ToCheckInst_LFInst_18_LFInst_0_n3,
         Red_ToCheckInst_LFInst_18_LFInst_1_n3,
         Red_ToCheckInst_LFInst_18_LFInst_2_n3,
         Red_ToCheckInst_LFInst_19_LFInst_0_n3,
         Red_ToCheckInst_LFInst_19_LFInst_1_n3,
         Red_ToCheckInst_LFInst_19_LFInst_2_n3,
         Red_ToCheckInst_LFInst_20_LFInst_0_n3,
         Red_ToCheckInst_LFInst_20_LFInst_1_n3,
         Red_ToCheckInst_LFInst_20_LFInst_2_n3,
         Red_ToCheckInst_LFInst_21_LFInst_0_n3,
         Red_ToCheckInst_LFInst_21_LFInst_1_n3,
         Red_ToCheckInst_LFInst_21_LFInst_2_n3,
         Red_ToCheckInst_LFInst_22_LFInst_0_n3,
         Red_ToCheckInst_LFInst_22_LFInst_1_n3,
         Red_ToCheckInst_LFInst_22_LFInst_2_n3,
         Red_ToCheckInst_LFInst_23_LFInst_0_n3,
         Red_ToCheckInst_LFInst_23_LFInst_1_n3,
         Red_ToCheckInst_LFInst_23_LFInst_2_n3,
         Red_ToCheckInst_LFInst_24_LFInst_0_n3,
         Red_ToCheckInst_LFInst_24_LFInst_1_n3,
         Red_ToCheckInst_LFInst_24_LFInst_2_n3,
         Red_ToCheckInst_LFInst_25_LFInst_0_n3,
         Red_ToCheckInst_LFInst_25_LFInst_1_n3,
         Red_ToCheckInst_LFInst_25_LFInst_2_n3,
         Red_ToCheckInst_LFInst_26_LFInst_0_n3,
         Red_ToCheckInst_LFInst_26_LFInst_1_n3,
         Red_ToCheckInst_LFInst_26_LFInst_2_n3,
         Red_ToCheckInst_LFInst_27_LFInst_0_n3,
         Red_ToCheckInst_LFInst_27_LFInst_1_n3,
         Red_ToCheckInst_LFInst_27_LFInst_2_n3,
         Red_ToCheckInst_LFInst_28_LFInst_0_n3,
         Red_ToCheckInst_LFInst_28_LFInst_1_n3,
         Red_ToCheckInst_LFInst_28_LFInst_2_n3,
         Red_ToCheckInst_LFInst_29_LFInst_0_n3,
         Red_ToCheckInst_LFInst_29_LFInst_1_n3,
         Red_ToCheckInst_LFInst_29_LFInst_2_n3,
         Red_ToCheckInst_LFInst_30_LFInst_0_n3,
         Red_ToCheckInst_LFInst_30_LFInst_1_n3,
         Red_ToCheckInst_LFInst_30_LFInst_2_n3,
         Red_ToCheckInst_LFInst_31_LFInst_0_n3,
         Red_ToCheckInst_LFInst_31_LFInst_1_n3,
         Red_ToCheckInst_LFInst_31_LFInst_2_n3,
         Red_ToCheckInst_LFInst_32_LFInst_0_n3,
         Red_ToCheckInst_LFInst_32_LFInst_1_n3,
         Red_ToCheckInst_LFInst_32_LFInst_2_n3,
         Red_ToCheckInst_LFInst_33_LFInst_0_n3,
         Red_ToCheckInst_LFInst_33_LFInst_1_n3,
         Red_ToCheckInst_LFInst_33_LFInst_2_n3,
         Red_ToCheckInst_LFInst_34_LFInst_0_n3,
         Red_ToCheckInst_LFInst_34_LFInst_1_n3,
         Red_ToCheckInst_LFInst_34_LFInst_2_n3,
         Red_ToCheckInst_LFInst_35_LFInst_0_n3,
         Red_ToCheckInst_LFInst_35_LFInst_1_n3,
         Red_ToCheckInst_LFInst_35_LFInst_2_n3,
         Red_ToCheckInst_LFInst_36_LFInst_0_n3,
         Red_ToCheckInst_LFInst_36_LFInst_1_n3,
         Red_ToCheckInst_LFInst_36_LFInst_2_n3,
         Red_ToCheckInst_LFInst_37_LFInst_0_n3,
         Red_ToCheckInst_LFInst_37_LFInst_1_n3,
         Red_ToCheckInst_LFInst_37_LFInst_2_n3,
         Red_ToCheckInst_LFInst_38_LFInst_0_n3,
         Red_ToCheckInst_LFInst_38_LFInst_1_n3,
         Red_ToCheckInst_LFInst_38_LFInst_2_n3,
         Red_ToCheckInst_LFInst_39_LFInst_0_n3,
         Red_ToCheckInst_LFInst_39_LFInst_1_n3,
         Red_ToCheckInst_LFInst_39_LFInst_2_n3,
         Red_ToCheckInst_LFInst_40_LFInst_0_n3,
         Red_ToCheckInst_LFInst_40_LFInst_1_n3,
         Red_ToCheckInst_LFInst_40_LFInst_2_n3,
         Red_ToCheckInst_LFInst_41_LFInst_0_n3,
         Red_ToCheckInst_LFInst_41_LFInst_1_n3,
         Red_ToCheckInst_LFInst_41_LFInst_2_n3,
         Red_ToCheckInst_LFInst_42_LFInst_0_n3,
         Red_ToCheckInst_LFInst_42_LFInst_1_n3,
         Red_ToCheckInst_LFInst_42_LFInst_2_n3,
         Red_ToCheckInst_LFInst_43_LFInst_0_n3,
         Red_ToCheckInst_LFInst_43_LFInst_1_n3,
         Red_ToCheckInst_LFInst_43_LFInst_2_n3,
         Red_ToCheckInst_LFInst_44_LFInst_0_n3,
         Red_ToCheckInst_LFInst_44_LFInst_1_n3,
         Red_ToCheckInst_LFInst_44_LFInst_2_n3,
         Red_ToCheckInst_LFInst_45_LFInst_0_n3,
         Red_ToCheckInst_LFInst_45_LFInst_1_n3,
         Red_ToCheckInst_LFInst_45_LFInst_2_n3,
         Red_ToCheckInst_LFInst_46_LFInst_0_n3,
         Red_ToCheckInst_LFInst_46_LFInst_1_n3,
         Red_ToCheckInst_LFInst_46_LFInst_2_n3,
         Red_ToCheckInst_LFInst_47_LFInst_0_n3,
         Red_ToCheckInst_LFInst_47_LFInst_1_n3,
         Red_ToCheckInst_LFInst_47_LFInst_2_n3, Check1_CheckInst_0_n94,
         Check1_CheckInst_0_n93, Check1_CheckInst_0_n92,
         Check1_CheckInst_0_n91, Check1_CheckInst_0_n90,
         Check1_CheckInst_0_n89, Check1_CheckInst_0_n88,
         Check1_CheckInst_0_n87, Check1_CheckInst_0_n86,
         Check1_CheckInst_0_n85, Check1_CheckInst_0_n84,
         Check1_CheckInst_0_n83, Check1_CheckInst_0_n82,
         Check1_CheckInst_0_n81, Check1_CheckInst_0_n80,
         Check1_CheckInst_0_n79, Check1_CheckInst_0_n78,
         Check1_CheckInst_0_n77, Check1_CheckInst_0_n76,
         Check1_CheckInst_0_n75, Check1_CheckInst_0_n74,
         Check1_CheckInst_0_n73, Check1_CheckInst_0_n72,
         Check1_CheckInst_0_n71, Check1_CheckInst_0_n70,
         Check1_CheckInst_0_n69, Check1_CheckInst_0_n68,
         Check1_CheckInst_0_n67, Check1_CheckInst_0_n66,
         Check1_CheckInst_0_n65, Check1_CheckInst_0_n64,
         Check1_CheckInst_0_n63, Check1_CheckInst_0_n62,
         Check1_CheckInst_0_n61, Check1_CheckInst_0_n60,
         Check1_CheckInst_0_n59, Check1_CheckInst_0_n58,
         Check1_CheckInst_0_n57, Check1_CheckInst_0_n56,
         Check1_CheckInst_0_n55, Check1_CheckInst_0_n54,
         Check1_CheckInst_0_n53, Check1_CheckInst_0_n52,
         Check1_CheckInst_0_n51, Check1_CheckInst_0_n50,
         Check1_CheckInst_0_n49, Check1_CheckInst_0_n48,
         Check1_CheckInst_0_n47, Check1_CheckInst_0_n46,
         Check1_CheckInst_0_n45, Check1_CheckInst_0_n44,
         Check1_CheckInst_0_n43, Check1_CheckInst_0_n42,
         Check1_CheckInst_0_n41, Check1_CheckInst_0_n40,
         Check1_CheckInst_0_n39, Check1_CheckInst_0_n38,
         Check1_CheckInst_0_n37, Check1_CheckInst_0_n36,
         Check1_CheckInst_0_n35, Check1_CheckInst_0_n34,
         Check1_CheckInst_0_n33, Check1_CheckInst_0_n32,
         Check1_CheckInst_0_n31, Check1_CheckInst_0_n30,
         Check1_CheckInst_0_n29, Check1_CheckInst_0_n28,
         Check1_CheckInst_0_n27, Check1_CheckInst_0_n26,
         Check1_CheckInst_0_n25, Check1_CheckInst_0_n24,
         Check1_CheckInst_0_n23, Check1_CheckInst_0_n22,
         Check1_CheckInst_0_n21, Check1_CheckInst_0_n20,
         Check1_CheckInst_0_n19, Check1_CheckInst_0_n18,
         Check1_CheckInst_0_n17, Check1_CheckInst_0_n16,
         Check1_CheckInst_0_n15, Check1_CheckInst_0_n14,
         Check1_CheckInst_0_n13, Check1_CheckInst_0_n12,
         Check1_CheckInst_0_n11, Check1_CheckInst_0_n10, Check1_CheckInst_0_n9,
         Check1_CheckInst_0_n8, Check1_CheckInst_0_n7, Check1_CheckInst_0_n6,
         Check1_CheckInst_0_n5, Check1_CheckInst_0_n4, Check1_CheckInst_0_n3,
         Check1_CheckInst_0_n2, Check1_CheckInst_0_n1, Check1_CheckInst_1_n96,
         Check1_CheckInst_1_n95, Check1_CheckInst_1_n94,
         Check1_CheckInst_1_n93, Check1_CheckInst_1_n92,
         Check1_CheckInst_1_n91, Check1_CheckInst_1_n90,
         Check1_CheckInst_1_n89, Check1_CheckInst_1_n88,
         Check1_CheckInst_1_n87, Check1_CheckInst_1_n86,
         Check1_CheckInst_1_n85, Check1_CheckInst_1_n84,
         Check1_CheckInst_1_n83, Check1_CheckInst_1_n82,
         Check1_CheckInst_1_n81, Check1_CheckInst_1_n80,
         Check1_CheckInst_1_n79, Check1_CheckInst_1_n78,
         Check1_CheckInst_1_n77, Check1_CheckInst_1_n76,
         Check1_CheckInst_1_n75, Check1_CheckInst_1_n74,
         Check1_CheckInst_1_n73, Check1_CheckInst_1_n72,
         Check1_CheckInst_1_n71, Check1_CheckInst_1_n70,
         Check1_CheckInst_1_n69, Check1_CheckInst_1_n68,
         Check1_CheckInst_1_n67, Check1_CheckInst_1_n66,
         Check1_CheckInst_1_n65, Check1_CheckInst_1_n64,
         Check1_CheckInst_1_n63, Check1_CheckInst_1_n62,
         Check1_CheckInst_1_n61, Check1_CheckInst_1_n60,
         Check1_CheckInst_1_n59, Check1_CheckInst_1_n58,
         Check1_CheckInst_1_n57, Check1_CheckInst_1_n56,
         Check1_CheckInst_1_n55, Check1_CheckInst_1_n54,
         Check1_CheckInst_1_n53, Check1_CheckInst_1_n52,
         Check1_CheckInst_1_n51, Check1_CheckInst_1_n50,
         Check1_CheckInst_1_n49, Check1_CheckInst_1_n48,
         Check1_CheckInst_1_n47, Check1_CheckInst_1_n46,
         Check1_CheckInst_1_n45, Check1_CheckInst_1_n44,
         Check1_CheckInst_1_n43, Check1_CheckInst_1_n42,
         Check1_CheckInst_1_n41, Check1_CheckInst_1_n40,
         Check1_CheckInst_1_n39, Check1_CheckInst_1_n38,
         Check1_CheckInst_1_n37, Check1_CheckInst_1_n36,
         Check1_CheckInst_1_n35, Check1_CheckInst_1_n34,
         Check1_CheckInst_1_n33, Check1_CheckInst_1_n32,
         Check1_CheckInst_1_n31, Check1_CheckInst_1_n30,
         Check1_CheckInst_1_n29, Check1_CheckInst_1_n28,
         Check1_CheckInst_1_n27, Check1_CheckInst_1_n26,
         Check1_CheckInst_1_n25, Check1_CheckInst_1_n24,
         Check1_CheckInst_1_n23, Check1_CheckInst_1_n22,
         Check1_CheckInst_1_n21, Check1_CheckInst_1_n20,
         Check1_CheckInst_1_n19, Check1_CheckInst_1_n18,
         Check1_CheckInst_1_n17, Check1_CheckInst_1_n16,
         Check1_CheckInst_1_n15, Check1_CheckInst_1_n14,
         Check1_CheckInst_1_n13, Check1_CheckInst_1_n12,
         Check1_CheckInst_1_n11, Check1_CheckInst_1_n10, Check1_CheckInst_1_n9,
         Check1_CheckInst_1_n8, Check1_CheckInst_1_n7, Check1_CheckInst_1_n6,
         Check1_CheckInst_1_n5, Check1_CheckInst_1_n4, Check1_CheckInst_1_n3,
         Check1_CheckInst_2_n96, Check1_CheckInst_2_n95,
         Check1_CheckInst_2_n94, Check1_CheckInst_2_n93,
         Check1_CheckInst_2_n92, Check1_CheckInst_2_n91,
         Check1_CheckInst_2_n90, Check1_CheckInst_2_n89,
         Check1_CheckInst_2_n88, Check1_CheckInst_2_n87,
         Check1_CheckInst_2_n86, Check1_CheckInst_2_n85,
         Check1_CheckInst_2_n84, Check1_CheckInst_2_n83,
         Check1_CheckInst_2_n82, Check1_CheckInst_2_n81,
         Check1_CheckInst_2_n80, Check1_CheckInst_2_n79,
         Check1_CheckInst_2_n78, Check1_CheckInst_2_n77,
         Check1_CheckInst_2_n76, Check1_CheckInst_2_n75,
         Check1_CheckInst_2_n74, Check1_CheckInst_2_n73,
         Check1_CheckInst_2_n72, Check1_CheckInst_2_n71,
         Check1_CheckInst_2_n70, Check1_CheckInst_2_n69,
         Check1_CheckInst_2_n68, Check1_CheckInst_2_n67,
         Check1_CheckInst_2_n66, Check1_CheckInst_2_n65,
         Check1_CheckInst_2_n64, Check1_CheckInst_2_n63,
         Check1_CheckInst_2_n62, Check1_CheckInst_2_n61,
         Check1_CheckInst_2_n60, Check1_CheckInst_2_n59,
         Check1_CheckInst_2_n58, Check1_CheckInst_2_n57,
         Check1_CheckInst_2_n56, Check1_CheckInst_2_n55,
         Check1_CheckInst_2_n54, Check1_CheckInst_2_n53,
         Check1_CheckInst_2_n52, Check1_CheckInst_2_n51,
         Check1_CheckInst_2_n50, Check1_CheckInst_2_n49,
         Check1_CheckInst_2_n48, Check1_CheckInst_2_n47,
         Check1_CheckInst_2_n46, Check1_CheckInst_2_n45,
         Check1_CheckInst_2_n44, Check1_CheckInst_2_n43,
         Check1_CheckInst_2_n42, Check1_CheckInst_2_n41,
         Check1_CheckInst_2_n40, Check1_CheckInst_2_n39,
         Check1_CheckInst_2_n38, Check1_CheckInst_2_n37,
         Check1_CheckInst_2_n36, Check1_CheckInst_2_n35,
         Check1_CheckInst_2_n34, Check1_CheckInst_2_n33,
         Check1_CheckInst_2_n32, Check1_CheckInst_2_n31,
         Check1_CheckInst_2_n30, Check1_CheckInst_2_n29,
         Check1_CheckInst_2_n28, Check1_CheckInst_2_n27,
         Check1_CheckInst_2_n26, Check1_CheckInst_2_n25,
         Check1_CheckInst_2_n24, Check1_CheckInst_2_n23,
         Check1_CheckInst_2_n22, Check1_CheckInst_2_n21,
         Check1_CheckInst_2_n20, Check1_CheckInst_2_n19,
         Check1_CheckInst_2_n18, Check1_CheckInst_2_n17,
         Check1_CheckInst_2_n16, Check1_CheckInst_2_n15,
         Check1_CheckInst_2_n14, Check1_CheckInst_2_n13,
         Check1_CheckInst_2_n12, Check1_CheckInst_2_n11,
         Check1_CheckInst_2_n10, Check1_CheckInst_2_n9, Check1_CheckInst_2_n8,
         Check1_CheckInst_2_n7, Check1_CheckInst_2_n6, Check1_CheckInst_2_n5,
         Check1_CheckInst_2_n4, Check1_CheckInst_2_n3;
  wire   [63:0] AddRoundKeyOutput;
  wire   [28:16] ShiftRowsOutput;
  wire   [47:0] Red_Plaintext;
  wire   [47:0] Red_RoundKey;
  wire   [47:0] Red_AddRoundKeyOutput;
  wire   [47:0] Red_ShiftRowsOutput;
  wire   [47:0] Red_MC_output;
  wire   [143:0] Red_SignaltoCheck;
  wire   [2:0] Error;
  wire   [3:0] MCInst_MC0_v3_3;
  wire   [3:0] MCInst_MC0_v3_2;
  wire   [3:0] MCInst_MC0_v3_1;
  wire   [3:1] MCInst_MC0_v3_0;
  wire   [3:0] MCInst_MC0_v2_3;
  wire   [3:0] MCInst_MC0_v2_2;
  wire   [3:0] MCInst_MC0_v2_1;
  wire   [3:1] MCInst_MC0_v2_0;
  wire   [3:1] MCInst_MC0_v1_3;
  wire   [3:0] MCInst_MC0_v1_2;
  wire   [3:0] MCInst_MC0_v1_1;
  wire   [3:1] MCInst_MC0_v0_3;
  wire   [3:0] MCInst_MC0_v0_2;
  wire   [3:1] MCInst_MC0_v0_1;
  wire   [2:1] MCInst_MC0_v0_0;
  wire   [3:0] MCInst_MC1_v3_3;
  wire   [3:0] MCInst_MC1_v3_2;
  wire   [3:0] MCInst_MC1_v3_1;
  wire   [3:1] MCInst_MC1_v3_0;
  wire   [3:0] MCInst_MC1_v2_3;
  wire   [3:0] MCInst_MC1_v2_2;
  wire   [3:0] MCInst_MC1_v2_1;
  wire   [3:1] MCInst_MC1_v2_0;
  wire   [3:1] MCInst_MC1_v1_3;
  wire   [3:0] MCInst_MC1_v1_2;
  wire   [3:0] MCInst_MC1_v1_1;
  wire   [3:1] MCInst_MC1_v0_3;
  wire   [3:0] MCInst_MC1_v0_2;
  wire   [3:1] MCInst_MC1_v0_1;
  wire   [2:1] MCInst_MC1_v0_0;
  wire   [3:0] MCInst_MC2_v3_3;
  wire   [3:0] MCInst_MC2_v3_2;
  wire   [3:0] MCInst_MC2_v3_1;
  wire   [3:1] MCInst_MC2_v3_0;
  wire   [3:0] MCInst_MC2_v2_3;
  wire   [3:0] MCInst_MC2_v2_2;
  wire   [3:0] MCInst_MC2_v2_1;
  wire   [3:1] MCInst_MC2_v2_0;
  wire   [3:1] MCInst_MC2_v1_3;
  wire   [3:0] MCInst_MC2_v1_2;
  wire   [3:0] MCInst_MC2_v1_1;
  wire   [3:1] MCInst_MC2_v0_3;
  wire   [3:0] MCInst_MC2_v0_2;
  wire   [3:1] MCInst_MC2_v0_1;
  wire   [2:1] MCInst_MC2_v0_0;
  wire   [3:0] MCInst_MC3_v3_3;
  wire   [3:0] MCInst_MC3_v3_2;
  wire   [3:0] MCInst_MC3_v3_1;
  wire   [3:1] MCInst_MC3_v3_0;
  wire   [3:0] MCInst_MC3_v2_3;
  wire   [3:0] MCInst_MC3_v2_2;
  wire   [3:0] MCInst_MC3_v2_1;
  wire   [3:1] MCInst_MC3_v2_0;
  wire   [3:1] MCInst_MC3_v1_3;
  wire   [3:0] MCInst_MC3_v1_2;
  wire   [3:0] MCInst_MC3_v1_1;
  wire   [3:1] MCInst_MC3_v0_3;
  wire   [3:0] MCInst_MC3_v0_2;
  wire   [3:1] MCInst_MC3_v0_1;
  wire   [2:1] MCInst_MC3_v0_0;
  wire   [2:0] Red_MCInst_MC0_v3_3;
  wire   [2:0] Red_MCInst_MC0_v3_2;
  wire   [2:1] Red_MCInst_MC0_v3_1;
  wire   [2:0] Red_MCInst_MC0_v3_0;
  wire   [2:0] Red_MCInst_MC0_v2_3;
  wire   [2:0] Red_MCInst_MC0_v2_2;
  wire   [2:0] Red_MCInst_MC0_v2_1;
  wire   [2:0] Red_MCInst_MC0_v2_0;
  wire   [2:0] Red_MCInst_MC0_v1_3;
  wire   [2:0] Red_MCInst_MC0_v1_2;
  wire   [2:1] Red_MCInst_MC0_v1_1;
  wire   [2:0] Red_MCInst_MC0_v1_0;
  wire   [2:0] Red_MCInst_MC0_v0_3;
  wire   [2:0] Red_MCInst_MC0_v0_2;
  wire   [2:0] Red_MCInst_MC0_v0_1;
  wire   [2:0] Red_MCInst_MC0_v0_0;
  wire   [2:0] Red_MCInst_MC1_v3_3;
  wire   [2:0] Red_MCInst_MC1_v3_2;
  wire   [2:1] Red_MCInst_MC1_v3_1;
  wire   [2:0] Red_MCInst_MC1_v3_0;
  wire   [2:0] Red_MCInst_MC1_v2_3;
  wire   [2:0] Red_MCInst_MC1_v2_2;
  wire   [2:0] Red_MCInst_MC1_v2_1;
  wire   [2:0] Red_MCInst_MC1_v2_0;
  wire   [2:0] Red_MCInst_MC1_v1_3;
  wire   [2:0] Red_MCInst_MC1_v1_2;
  wire   [2:1] Red_MCInst_MC1_v1_1;
  wire   [2:0] Red_MCInst_MC1_v1_0;
  wire   [2:0] Red_MCInst_MC1_v0_3;
  wire   [2:0] Red_MCInst_MC1_v0_2;
  wire   [2:0] Red_MCInst_MC1_v0_1;
  wire   [2:0] Red_MCInst_MC1_v0_0;
  wire   [2:0] Red_MCInst_MC2_v3_3;
  wire   [2:0] Red_MCInst_MC2_v3_2;
  wire   [2:1] Red_MCInst_MC2_v3_1;
  wire   [2:0] Red_MCInst_MC2_v3_0;
  wire   [2:0] Red_MCInst_MC2_v2_3;
  wire   [2:0] Red_MCInst_MC2_v2_2;
  wire   [2:0] Red_MCInst_MC2_v2_1;
  wire   [2:0] Red_MCInst_MC2_v2_0;
  wire   [2:0] Red_MCInst_MC2_v1_3;
  wire   [2:0] Red_MCInst_MC2_v1_2;
  wire   [2:1] Red_MCInst_MC2_v1_1;
  wire   [2:0] Red_MCInst_MC2_v1_0;
  wire   [2:0] Red_MCInst_MC2_v0_3;
  wire   [2:0] Red_MCInst_MC2_v0_2;
  wire   [2:0] Red_MCInst_MC2_v0_1;
  wire   [2:0] Red_MCInst_MC2_v0_0;
  wire   [2:0] Red_MCInst_MC3_v3_3;
  wire   [2:0] Red_MCInst_MC3_v3_2;
  wire   [2:1] Red_MCInst_MC3_v3_1;
  wire   [2:0] Red_MCInst_MC3_v3_0;
  wire   [2:0] Red_MCInst_MC3_v2_3;
  wire   [2:0] Red_MCInst_MC3_v2_2;
  wire   [2:0] Red_MCInst_MC3_v2_1;
  wire   [2:0] Red_MCInst_MC3_v2_0;
  wire   [2:0] Red_MCInst_MC3_v1_3;
  wire   [2:0] Red_MCInst_MC3_v1_2;
  wire   [2:1] Red_MCInst_MC3_v1_1;
  wire   [2:0] Red_MCInst_MC3_v1_0;
  wire   [2:0] Red_MCInst_MC3_v0_3;
  wire   [2:0] Red_MCInst_MC3_v0_2;
  wire   [2:0] Red_MCInst_MC3_v0_1;
  wire   [2:0] Red_MCInst_MC3_v0_0;

  AND2_X1 U6 ( .A1(Error[1]), .A2(Error[2]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(Error[0]), .A2(n4), .ZN(ErrorFlag) );
  XOR2_X2 AddKeyXOR_XORInst_0_0_U1 ( .A(Plaintext[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X2 AddKeyXOR_XORInst_0_1_U1 ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X2 AddKeyXOR_XORInst_0_2_U1 ( .A(Plaintext[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X2 AddKeyXOR_XORInst_0_3_U1 ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X2 AddKeyXOR_XORInst_1_0_U1 ( .A(Plaintext[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X2 AddKeyXOR_XORInst_1_1_U1 ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X2 AddKeyXOR_XORInst_1_2_U1 ( .A(Plaintext[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X2 AddKeyXOR_XORInst_1_3_U1 ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X2 AddKeyXOR_XORInst_2_0_U1 ( .A(Plaintext[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X2 AddKeyXOR_XORInst_2_1_U1 ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X2 AddKeyXOR_XORInst_2_2_U1 ( .A(Plaintext[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X2 AddKeyXOR_XORInst_2_3_U1 ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X2 AddKeyXOR_XORInst_3_0_U1 ( .A(Plaintext[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X2 AddKeyXOR_XORInst_3_1_U1 ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X2 AddKeyXOR_XORInst_3_2_U1 ( .A(Plaintext[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X2 AddKeyXOR_XORInst_3_3_U1 ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X2 AddKeyXOR_XORInst_4_0_U1 ( .A(Plaintext[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X2 AddKeyXOR_XORInst_4_1_U1 ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X2 AddKeyXOR_XORInst_4_2_U1 ( .A(Plaintext[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X2 AddKeyXOR_XORInst_4_3_U1 ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X2 AddKeyXOR_XORInst_5_0_U1 ( .A(Plaintext[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X2 AddKeyXOR_XORInst_5_1_U1 ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X2 AddKeyXOR_XORInst_5_2_U1 ( .A(Plaintext[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X2 AddKeyXOR_XORInst_5_3_U1 ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X2 AddKeyXOR_XORInst_6_0_U1 ( .A(Plaintext[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X2 AddKeyXOR_XORInst_6_1_U1 ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X2 AddKeyXOR_XORInst_6_2_U1 ( .A(Plaintext[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X2 AddKeyXOR_XORInst_6_3_U1 ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X2 AddKeyXOR_XORInst_7_0_U1 ( .A(Plaintext[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X2 AddKeyXOR_XORInst_7_1_U1 ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X2 AddKeyXOR_XORInst_7_2_U1 ( .A(Plaintext[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X2 AddKeyXOR_XORInst_7_3_U1 ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X2 AddKeyXOR_XORInst_8_0_U1 ( .A(Plaintext[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X2 AddKeyXOR_XORInst_8_1_U1 ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X2 AddKeyXOR_XORInst_8_2_U1 ( .A(Plaintext[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X2 AddKeyXOR_XORInst_8_3_U1 ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X2 AddKeyXOR_XORInst_9_0_U1 ( .A(Plaintext[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X2 AddKeyXOR_XORInst_9_1_U1 ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X2 AddKeyXOR_XORInst_9_2_U1 ( .A(Plaintext[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X2 AddKeyXOR_XORInst_9_3_U1 ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  XOR2_X2 AddKeyXOR_XORInst_10_0_U1 ( .A(Plaintext[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X2 AddKeyXOR_XORInst_10_1_U1 ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X2 AddKeyXOR_XORInst_10_2_U1 ( .A(Plaintext[42]), .B(Key[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X2 AddKeyXOR_XORInst_10_3_U1 ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X2 AddKeyXOR_XORInst_11_0_U1 ( .A(Plaintext[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X2 AddKeyXOR_XORInst_11_1_U1 ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X2 AddKeyXOR_XORInst_11_2_U1 ( .A(Plaintext[46]), .B(Key[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X2 AddKeyXOR_XORInst_11_3_U1 ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X2 AddKeyXOR_XORInst_12_0_U1 ( .A(Plaintext[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X2 AddKeyXOR_XORInst_12_1_U1 ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X2 AddKeyXOR_XORInst_12_2_U1 ( .A(Plaintext[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X2 AddKeyXOR_XORInst_12_3_U1 ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X2 AddKeyXOR_XORInst_13_0_U1 ( .A(Plaintext[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X2 AddKeyXOR_XORInst_13_1_U1 ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X2 AddKeyXOR_XORInst_13_2_U1 ( .A(Plaintext[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X2 AddKeyXOR_XORInst_13_3_U1 ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X2 AddKeyXOR_XORInst_14_0_U1 ( .A(Plaintext[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X2 AddKeyXOR_XORInst_14_1_U1 ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X2 AddKeyXOR_XORInst_14_2_U1 ( .A(Plaintext[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X2 AddKeyXOR_XORInst_14_3_U1 ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X2 AddKeyXOR_XORInst_15_0_U1 ( .A(Plaintext[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X2 AddKeyXOR_XORInst_15_1_U1 ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X2 AddKeyXOR_XORInst_15_2_U1 ( .A(Plaintext[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X2 AddKeyXOR_XORInst_15_3_U1 ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_0_U5 ( .A1(AddRoundKeyOutput[2]), .A2(
        SubCellInst_LFInst_0_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U4 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U3 ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_0_LFInst_0_n10), .ZN(MCInst_MC0_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_0_LFInst_0_n9), .B(SubCellInst_LFInst_0_LFInst_0_n8), .Z(SubCellInst_LFInst_0_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n24), .A2(
        SubCellInst_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U9 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U8 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n21), .A2(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n20), .A2(
        SubCellInst_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U5 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n19), .A2(
        SubCellInst_LFInst_0_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U3 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U2 ( .A(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_0_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n26), .A2(
        SubCellInst_LFInst_0_LFInst_1_n25), .ZN(Red_MCInst_MC0_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n25), .A2(
        SubCellInst_LFInst_0_LFInst_2_n28), .ZN(MCInst_MC0_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U7 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_0_LFInst_2_n26), .B(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n22), .A2(
        SubCellInst_LFInst_0_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_2_U3 ( .A(AddRoundKeyOutput[2]), .B(
        SubCellInst_LFInst_0_LFInst_2_n23), .Z(
        SubCellInst_LFInst_0_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U9 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n23), .A2(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U7 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n23), .A2(
        SubCellInst_LFInst_0_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n20), .A2(
        SubCellInst_LFInst_0_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4 ( .A1(AddRoundKeyOutput[2]), .A2(
        AddRoundKeyOutput[0]), .ZN(SubCellInst_LFInst_0_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_0_LFInst_3_U3 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n26), .A2(
        SubCellInst_LFInst_0_LFInst_3_n25), .ZN(Red_MCInst_MC0_v3_1[2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_0_U5 ( .A1(AddRoundKeyOutput[6]), .A2(
        SubCellInst_LFInst_1_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U4 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U3 ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_1_LFInst_0_n10), .ZN(MCInst_MC3_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_1_LFInst_0_n9), .B(SubCellInst_LFInst_1_LFInst_0_n8), .Z(SubCellInst_LFInst_1_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n24), .A2(
        SubCellInst_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U9 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U8 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n21), .A2(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n20), .A2(
        SubCellInst_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U5 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n19), .A2(
        SubCellInst_LFInst_1_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U3 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U2 ( .A(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_1_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n26), .A2(
        SubCellInst_LFInst_1_LFInst_1_n25), .ZN(Red_MCInst_MC3_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n25), .A2(
        SubCellInst_LFInst_1_LFInst_2_n28), .ZN(MCInst_MC3_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U7 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_1_LFInst_2_n26), .B(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n22), .A2(
        SubCellInst_LFInst_1_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_2_U3 ( .A(AddRoundKeyOutput[6]), .B(
        SubCellInst_LFInst_1_LFInst_2_n23), .Z(
        SubCellInst_LFInst_1_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U2 ( .A1(AddRoundKeyOutput[5]), .A2(
        AddRoundKeyOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U9 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n23), .A2(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U7 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n23), .A2(
        SubCellInst_LFInst_1_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n20), .A2(
        SubCellInst_LFInst_1_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4 ( .A1(AddRoundKeyOutput[6]), .A2(
        AddRoundKeyOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_1_LFInst_3_U3 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U2 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n26), .A2(
        SubCellInst_LFInst_1_LFInst_3_n25), .ZN(Red_MCInst_MC3_v3_1[2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_0_U5 ( .A1(AddRoundKeyOutput[10]), .A2(
        SubCellInst_LFInst_2_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U4 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U3 ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .Z(SubCellInst_LFInst_2_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_2_LFInst_0_n10), .ZN(MCInst_MC2_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_2_LFInst_0_n9), .B(SubCellInst_LFInst_2_LFInst_0_n8), .Z(SubCellInst_LFInst_2_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n24), .A2(
        SubCellInst_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U9 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U8 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n21), .A2(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n20), .A2(
        SubCellInst_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U5 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n19), .A2(
        SubCellInst_LFInst_2_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U3 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U2 ( .A(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_2_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n26), .A2(
        SubCellInst_LFInst_2_LFInst_1_n25), .ZN(Red_MCInst_MC2_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n25), .A2(
        SubCellInst_LFInst_2_LFInst_2_n28), .ZN(MCInst_MC2_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U7 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_2_LFInst_2_n26), .B(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n22), .A2(
        SubCellInst_LFInst_2_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_2_U3 ( .A(AddRoundKeyOutput[10]), .B(
        SubCellInst_LFInst_2_LFInst_2_n23), .Z(
        SubCellInst_LFInst_2_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U2 ( .A1(AddRoundKeyOutput[9]), .A2(
        AddRoundKeyOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U1 ( .A(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U9 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n23), .A2(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U7 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n23), .A2(
        SubCellInst_LFInst_2_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n20), .A2(
        SubCellInst_LFInst_2_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4 ( .A1(AddRoundKeyOutput[10]), .A2(
        AddRoundKeyOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_2_LFInst_3_U3 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U2 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n26), .A2(
        SubCellInst_LFInst_2_LFInst_3_n25), .ZN(Red_MCInst_MC2_v3_1[2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_0_U5 ( .A1(AddRoundKeyOutput[14]), .A2(
        SubCellInst_LFInst_3_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U4 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U3 ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .Z(SubCellInst_LFInst_3_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_3_LFInst_0_n10), .ZN(MCInst_MC1_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_3_LFInst_0_n9), .B(SubCellInst_LFInst_3_LFInst_0_n8), .Z(SubCellInst_LFInst_3_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n24), .A2(
        SubCellInst_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U9 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U8 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n21), .A2(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n20), .A2(
        SubCellInst_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U5 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n19), .A2(
        SubCellInst_LFInst_3_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U3 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U2 ( .A(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_3_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n26), .A2(
        SubCellInst_LFInst_3_LFInst_1_n25), .ZN(Red_MCInst_MC1_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n25), .A2(
        SubCellInst_LFInst_3_LFInst_2_n28), .ZN(MCInst_MC1_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U7 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_3_LFInst_2_n26), .B(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n22), .A2(
        SubCellInst_LFInst_3_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_2_U3 ( .A(AddRoundKeyOutput[14]), .B(
        SubCellInst_LFInst_3_LFInst_2_n23), .Z(
        SubCellInst_LFInst_3_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U2 ( .A1(AddRoundKeyOutput[13]), .A2(
        AddRoundKeyOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U1 ( .A(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U9 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n23), .A2(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U7 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n23), .A2(
        SubCellInst_LFInst_3_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n20), .A2(
        SubCellInst_LFInst_3_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4 ( .A1(AddRoundKeyOutput[14]), .A2(
        AddRoundKeyOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_3_LFInst_3_U3 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U2 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n26), .A2(
        SubCellInst_LFInst_3_LFInst_3_n25), .ZN(Red_MCInst_MC1_v3_1[2]) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_4_LFInst_0_n8), .B(SubCellInst_LFInst_4_LFInst_0_n7), .ZN(ShiftRowsOutput[24]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(AddRoundKeyOutput[18]), .A2(
        SubCellInst_LFInst_4_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U2 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n24), .A2(
        SubCellInst_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U9 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U8 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n21), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n20), .A2(
        SubCellInst_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U5 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n19), .A2(
        SubCellInst_LFInst_4_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U3 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U2 ( .A(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n26), .A2(
        SubCellInst_LFInst_4_LFInst_1_n25), .ZN(MCInst_MC1_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U9 ( .A1(AddRoundKeyOutput[18]), .A2(
        SubCellInst_LFInst_4_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_2_U8 ( .A1(AddRoundKeyOutput[17]), .A2(
        SubCellInst_LFInst_4_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U7 ( .A(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n25), .A2(
        SubCellInst_LFInst_4_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_4_LFInst_2_n23), .B(AddRoundKeyOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n22), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_2_U2 ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_4_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n29), .A2(
        SubCellInst_LFInst_4_LFInst_2_n28), .ZN(MCInst_MC1_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n25), .A2(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n25), .A2(
        SubCellInst_LFInst_4_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n22), .A2(
        SubCellInst_LFInst_4_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U6 ( .A1(AddRoundKeyOutput[18]), .A2(
        AddRoundKeyOutput[16]), .ZN(SubCellInst_LFInst_4_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_4_LFInst_3_U5 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_3_U3 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U2 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_4_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n19), .A2(
        SubCellInst_LFInst_4_LFInst_3_n20), .ZN(Red_MCInst_MC1_v2_2[1]) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_5_LFInst_0_n8), .B(SubCellInst_LFInst_5_LFInst_0_n7), .ZN(ShiftRowsOutput[28]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(AddRoundKeyOutput[22]), .A2(
        SubCellInst_LFInst_5_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U2 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n24), .A2(
        SubCellInst_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U9 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U8 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n21), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n20), .A2(
        SubCellInst_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U5 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n19), .A2(
        SubCellInst_LFInst_5_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U3 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U2 ( .A(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n26), .A2(
        SubCellInst_LFInst_5_LFInst_1_n25), .ZN(MCInst_MC0_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U9 ( .A1(AddRoundKeyOutput[22]), .A2(
        SubCellInst_LFInst_5_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_2_U8 ( .A1(AddRoundKeyOutput[21]), .A2(
        SubCellInst_LFInst_5_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U7 ( .A(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n25), .A2(
        SubCellInst_LFInst_5_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_5_LFInst_2_n23), .B(AddRoundKeyOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n22), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_2_U2 ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_5_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n29), .A2(
        SubCellInst_LFInst_5_LFInst_2_n28), .ZN(MCInst_MC0_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n25), .A2(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n25), .A2(
        SubCellInst_LFInst_5_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n22), .A2(
        SubCellInst_LFInst_5_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U6 ( .A1(AddRoundKeyOutput[22]), .A2(
        AddRoundKeyOutput[20]), .ZN(SubCellInst_LFInst_5_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_5_LFInst_3_U5 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_3_U3 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U2 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_5_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n19), .A2(
        SubCellInst_LFInst_5_LFInst_3_n20), .ZN(Red_MCInst_MC0_v2_2[1]) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_6_LFInst_0_n8), .B(SubCellInst_LFInst_6_LFInst_0_n7), .ZN(ShiftRowsOutput[16]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(AddRoundKeyOutput[26]), .A2(
        SubCellInst_LFInst_6_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U2 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .Z(SubCellInst_LFInst_6_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n24), .A2(
        SubCellInst_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U9 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U8 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n21), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n20), .A2(
        SubCellInst_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U5 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n19), .A2(
        SubCellInst_LFInst_6_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U3 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U2 ( .A(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n26), .A2(
        SubCellInst_LFInst_6_LFInst_1_n25), .ZN(MCInst_MC3_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U9 ( .A1(AddRoundKeyOutput[26]), .A2(
        SubCellInst_LFInst_6_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_2_U8 ( .A1(AddRoundKeyOutput[25]), .A2(
        SubCellInst_LFInst_6_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U7 ( .A(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n25), .A2(
        SubCellInst_LFInst_6_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_6_LFInst_2_n23), .B(AddRoundKeyOutput[26]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n22), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_2_U2 ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_6_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n29), .A2(
        SubCellInst_LFInst_6_LFInst_2_n28), .ZN(MCInst_MC3_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n25), .A2(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n25), .A2(
        SubCellInst_LFInst_6_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n22), .A2(
        SubCellInst_LFInst_6_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U6 ( .A1(AddRoundKeyOutput[26]), .A2(
        AddRoundKeyOutput[24]), .ZN(SubCellInst_LFInst_6_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_6_LFInst_3_U5 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_3_U3 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U2 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_6_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n19), .A2(
        SubCellInst_LFInst_6_LFInst_3_n20), .ZN(Red_MCInst_MC3_v2_2[1]) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_7_LFInst_0_n8), .B(SubCellInst_LFInst_7_LFInst_0_n7), .ZN(ShiftRowsOutput[20]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(AddRoundKeyOutput[30]), .A2(
        SubCellInst_LFInst_7_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U2 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .Z(SubCellInst_LFInst_7_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n24), .A2(
        SubCellInst_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U9 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U8 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n21), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n20), .A2(
        SubCellInst_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U5 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n19), .A2(
        SubCellInst_LFInst_7_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U3 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U2 ( .A(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n26), .A2(
        SubCellInst_LFInst_7_LFInst_1_n25), .ZN(MCInst_MC2_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U9 ( .A1(AddRoundKeyOutput[30]), .A2(
        SubCellInst_LFInst_7_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_2_U8 ( .A1(AddRoundKeyOutput[29]), .A2(
        SubCellInst_LFInst_7_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U7 ( .A(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n25), .A2(
        SubCellInst_LFInst_7_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_7_LFInst_2_n23), .B(AddRoundKeyOutput[30]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n22), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_2_U2 ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_7_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n29), .A2(
        SubCellInst_LFInst_7_LFInst_2_n28), .ZN(MCInst_MC2_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n25), .A2(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n25), .A2(
        SubCellInst_LFInst_7_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n22), .A2(
        SubCellInst_LFInst_7_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U6 ( .A1(AddRoundKeyOutput[30]), .A2(
        AddRoundKeyOutput[28]), .ZN(SubCellInst_LFInst_7_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_7_LFInst_3_U5 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_3_U3 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U2 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_7_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n19), .A2(
        SubCellInst_LFInst_7_LFInst_3_n20), .ZN(Red_MCInst_MC2_v2_2[1]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_0_U5 ( .A1(AddRoundKeyOutput[34]), .A2(
        SubCellInst_LFInst_8_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U4 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U3 ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_8_LFInst_0_n12), .ZN(MCInst_MC2_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_8_LFInst_0_n11), .B(
        SubCellInst_LFInst_8_LFInst_0_n10), .Z(
        SubCellInst_LFInst_8_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n26), .A2(
        SubCellInst_LFInst_8_LFInst_1_n25), .ZN(MCInst_MC2_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n24), .A2(
        SubCellInst_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U8 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U7 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n21), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n20), .A2(
        SubCellInst_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n19), .A2(
        SubCellInst_LFInst_8_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U1 ( .A(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n24), .A2(
        SubCellInst_LFInst_8_LFInst_2_n28), .ZN(MCInst_MC2_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U7 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n26), .A2(
        SubCellInst_LFInst_8_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n28) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U6 ( .A(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n27) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_8_LFInst_2_n25), .B(AddRoundKeyOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n25) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n23), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n24) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U2 ( .A(
        SubCellInst_LFInst_8_LFInst_2_n22), .B(AddRoundKeyOutput[33]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n23) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_2_U1 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U9 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n23), .A2(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U7 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n23), .A2(
        SubCellInst_LFInst_8_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n20), .A2(
        SubCellInst_LFInst_8_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U4 ( .A1(AddRoundKeyOutput[34]), .A2(
        AddRoundKeyOutput[32]), .ZN(SubCellInst_LFInst_8_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_8_LFInst_3_U3 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U2 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n26), .A2(
        SubCellInst_LFInst_8_LFInst_3_n25), .ZN(Red_MCInst_MC2_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_0_U5 ( .A1(AddRoundKeyOutput[38]), .A2(
        SubCellInst_LFInst_9_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U4 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U3 ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_9_LFInst_0_n12), .ZN(MCInst_MC1_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_9_LFInst_0_n11), .B(
        SubCellInst_LFInst_9_LFInst_0_n10), .Z(
        SubCellInst_LFInst_9_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n26), .A2(
        SubCellInst_LFInst_9_LFInst_1_n25), .ZN(MCInst_MC1_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n24), .A2(
        SubCellInst_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U8 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U7 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n21), .A2(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n20), .A2(
        SubCellInst_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n19), .A2(
        SubCellInst_LFInst_9_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U1 ( .A(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n25), .A2(
        SubCellInst_LFInst_9_LFInst_2_n28), .ZN(MCInst_MC1_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U7 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_9_LFInst_2_n26), .B(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n22), .A2(
        SubCellInst_LFInst_9_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_2_U3 ( .A(AddRoundKeyOutput[38]), .B(
        SubCellInst_LFInst_9_LFInst_2_n23), .Z(
        SubCellInst_LFInst_9_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U2 ( .A1(AddRoundKeyOutput[37]), .A2(
        AddRoundKeyOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U1 ( .A(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U9 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n23), .A2(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U7 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n23), .A2(
        SubCellInst_LFInst_9_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n20), .A2(
        SubCellInst_LFInst_9_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U4 ( .A1(AddRoundKeyOutput[38]), .A2(
        AddRoundKeyOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_9_LFInst_3_U3 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U2 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n26), .A2(
        SubCellInst_LFInst_9_LFInst_3_n25), .ZN(Red_MCInst_MC1_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_0_U5 ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U4 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U3 ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .Z(SubCellInst_LFInst_10_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_10_LFInst_0_n12), .ZN(MCInst_MC0_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_10_LFInst_0_n11), .B(
        SubCellInst_LFInst_10_LFInst_0_n10), .Z(
        SubCellInst_LFInst_10_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n26), .A2(
        SubCellInst_LFInst_10_LFInst_1_n25), .ZN(MCInst_MC0_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n24), .A2(
        SubCellInst_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U8 ( .A1(AddRoundKeyOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U7 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n21), .A2(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n20), .A2(
        SubCellInst_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n19), .A2(
        SubCellInst_LFInst_10_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U1 ( .A(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n25), .A2(
        SubCellInst_LFInst_10_LFInst_2_n28), .ZN(MCInst_MC0_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U7 ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_10_LFInst_2_n26), .B(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(AddRoundKeyOutput[40]), .A2(
        AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n22), .A2(
        SubCellInst_LFInst_10_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_2_U3 ( .A(AddRoundKeyOutput[42]), .B(
        SubCellInst_LFInst_10_LFInst_2_n23), .Z(
        SubCellInst_LFInst_10_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U2 ( .A1(AddRoundKeyOutput[41]), 
        .A2(AddRoundKeyOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U1 ( .A(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U9 ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n23), .A2(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U7 ( .A1(AddRoundKeyOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n23), .A2(
        SubCellInst_LFInst_10_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n20), .A2(
        SubCellInst_LFInst_10_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U4 ( .A1(AddRoundKeyOutput[42]), .A2(
        AddRoundKeyOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_10_LFInst_3_U3 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U2 ( .A1(AddRoundKeyOutput[40]), .A2(
        AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n26), .A2(
        SubCellInst_LFInst_10_LFInst_3_n25), .ZN(Red_MCInst_MC0_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_0_U5 ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U4 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U3 ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .Z(SubCellInst_LFInst_11_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_11_LFInst_0_n12), .ZN(MCInst_MC3_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_11_LFInst_0_n11), .B(
        SubCellInst_LFInst_11_LFInst_0_n10), .Z(
        SubCellInst_LFInst_11_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n26), .A2(
        SubCellInst_LFInst_11_LFInst_1_n25), .ZN(MCInst_MC3_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U9 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n24), .A2(
        SubCellInst_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U8 ( .A1(AddRoundKeyOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U7 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n21), .A2(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U5 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n20), .A2(
        SubCellInst_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U3 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n19), .A2(
        SubCellInst_LFInst_11_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U1 ( .A(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n25), .A2(
        SubCellInst_LFInst_11_LFInst_2_n28), .ZN(MCInst_MC3_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U7 ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_11_LFInst_2_n26), .B(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(AddRoundKeyOutput[44]), .A2(
        AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n22), .A2(
        SubCellInst_LFInst_11_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_2_U3 ( .A(AddRoundKeyOutput[46]), .B(
        SubCellInst_LFInst_11_LFInst_2_n23), .Z(
        SubCellInst_LFInst_11_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U2 ( .A1(AddRoundKeyOutput[45]), 
        .A2(AddRoundKeyOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U9 ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n23), .A2(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U7 ( .A1(AddRoundKeyOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n23), .A2(
        SubCellInst_LFInst_11_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n20), .A2(
        SubCellInst_LFInst_11_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U4 ( .A1(AddRoundKeyOutput[46]), .A2(
        AddRoundKeyOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_11_LFInst_3_U3 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U2 ( .A1(AddRoundKeyOutput[44]), .A2(
        AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n26), .A2(
        SubCellInst_LFInst_11_LFInst_3_n25), .ZN(Red_MCInst_MC3_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_0_U5 ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U4 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U3 ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_12_LFInst_0_n9), .ZN(Red_MCInst_MC3_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_12_LFInst_0_n8), .B(
        SubCellInst_LFInst_12_LFInst_0_n7), .Z(
        SubCellInst_LFInst_12_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n24), .A2(
        SubCellInst_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U9 ( .A1(AddRoundKeyOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U8 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n21), .A2(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n20), .A2(
        SubCellInst_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U5 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n19), .A2(
        SubCellInst_LFInst_12_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U3 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U2 ( .A(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n26), .A2(
        SubCellInst_LFInst_12_LFInst_1_n25), .ZN(Red_MCInst_MC3_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n24), .A2(
        SubCellInst_LFInst_12_LFInst_2_n28), .ZN(MCInst_MC3_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U7 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n26), .A2(
        SubCellInst_LFInst_12_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n28) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U6 ( .A(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n27) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_12_LFInst_2_n25), .B(AddRoundKeyOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n25) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n23), .A2(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n24) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U2 ( .A(
        SubCellInst_LFInst_12_LFInst_2_n22), .B(AddRoundKeyOutput[49]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n23) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_2_U1 ( .A1(AddRoundKeyOutput[48]), .A2(
        AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U9 ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n23), .A2(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U7 ( .A1(AddRoundKeyOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n23), .A2(
        SubCellInst_LFInst_12_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n20), .A2(
        SubCellInst_LFInst_12_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U4 ( .A1(AddRoundKeyOutput[50]), .A2(
        AddRoundKeyOutput[48]), .ZN(SubCellInst_LFInst_12_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_12_LFInst_3_U3 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U2 ( .A1(AddRoundKeyOutput[48]), .A2(
        AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n26), .A2(
        SubCellInst_LFInst_12_LFInst_3_n25), .ZN(Red_MCInst_MC3_v0_1[0]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_0_U5 ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U4 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U3 ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_13_LFInst_0_n9), .ZN(Red_MCInst_MC2_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_13_LFInst_0_n8), .B(
        SubCellInst_LFInst_13_LFInst_0_n7), .Z(
        SubCellInst_LFInst_13_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n24), .A2(
        SubCellInst_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U9 ( .A1(AddRoundKeyOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U8 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n21), .A2(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n20), .A2(
        SubCellInst_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U5 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n19), .A2(
        SubCellInst_LFInst_13_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U2 ( .A(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n26), .A2(
        SubCellInst_LFInst_13_LFInst_1_n25), .ZN(Red_MCInst_MC2_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U9 ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_2_U8 ( .A1(AddRoundKeyOutput[53]), .A2(
        SubCellInst_LFInst_13_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U7 ( .A(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n25), .A2(
        SubCellInst_LFInst_13_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_13_LFInst_2_n23), .B(AddRoundKeyOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n22), .A2(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_2_U2 ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n29), .A2(
        SubCellInst_LFInst_13_LFInst_2_n28), .ZN(MCInst_MC2_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U9 ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n23), .A2(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U7 ( .A1(AddRoundKeyOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n23), .A2(
        SubCellInst_LFInst_13_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n20), .A2(
        SubCellInst_LFInst_13_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U4 ( .A1(AddRoundKeyOutput[54]), .A2(
        AddRoundKeyOutput[52]), .ZN(SubCellInst_LFInst_13_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_13_LFInst_3_U3 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U2 ( .A1(AddRoundKeyOutput[52]), .A2(
        AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n26), .A2(
        SubCellInst_LFInst_13_LFInst_3_n25), .ZN(Red_MCInst_MC2_v0_1[0]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_0_U5 ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U4 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U3 ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .Z(SubCellInst_LFInst_14_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_14_LFInst_0_n9), .ZN(Red_MCInst_MC1_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_14_LFInst_0_n8), .B(
        SubCellInst_LFInst_14_LFInst_0_n7), .Z(
        SubCellInst_LFInst_14_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n24), .A2(
        SubCellInst_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U9 ( .A1(AddRoundKeyOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U8 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n21), .A2(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n20), .A2(
        SubCellInst_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U5 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n19), .A2(
        SubCellInst_LFInst_14_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U3 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U2 ( .A(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n26), .A2(
        SubCellInst_LFInst_14_LFInst_1_n25), .ZN(Red_MCInst_MC1_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n24), .A2(
        SubCellInst_LFInst_14_LFInst_2_n28), .ZN(MCInst_MC1_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U7 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n26), .A2(
        SubCellInst_LFInst_14_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n28) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U6 ( .A(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n27) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_14_LFInst_2_n25), .B(AddRoundKeyOutput[58]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n25) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n23), .A2(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n24) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U2 ( .A(
        SubCellInst_LFInst_14_LFInst_2_n22), .B(AddRoundKeyOutput[57]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n23) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_2_U1 ( .A1(AddRoundKeyOutput[56]), .A2(
        AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U9 ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n23), .A2(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U7 ( .A1(AddRoundKeyOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n23), .A2(
        SubCellInst_LFInst_14_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n20), .A2(
        SubCellInst_LFInst_14_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U4 ( .A1(AddRoundKeyOutput[58]), .A2(
        AddRoundKeyOutput[56]), .ZN(SubCellInst_LFInst_14_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_14_LFInst_3_U3 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U2 ( .A1(AddRoundKeyOutput[56]), .A2(
        AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n26), .A2(
        SubCellInst_LFInst_14_LFInst_3_n25), .ZN(Red_MCInst_MC1_v0_1[0]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_0_U5 ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U4 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U3 ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .Z(SubCellInst_LFInst_15_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_15_LFInst_0_n9), .ZN(Red_MCInst_MC0_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_15_LFInst_0_n8), .B(
        SubCellInst_LFInst_15_LFInst_0_n7), .Z(
        SubCellInst_LFInst_15_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n24), .A2(
        SubCellInst_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U9 ( .A1(AddRoundKeyOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U8 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n21), .A2(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n20), .A2(
        SubCellInst_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U5 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n19), .A2(
        SubCellInst_LFInst_15_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U3 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U2 ( .A(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n26), .A2(
        SubCellInst_LFInst_15_LFInst_1_n25), .ZN(Red_MCInst_MC0_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n24), .A2(
        SubCellInst_LFInst_15_LFInst_2_n28), .ZN(MCInst_MC0_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U7 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n26), .A2(
        SubCellInst_LFInst_15_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n28) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U6 ( .A(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n27) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_15_LFInst_2_n25), .B(AddRoundKeyOutput[62]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n25) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n23), .A2(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n24) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U2 ( .A(
        SubCellInst_LFInst_15_LFInst_2_n22), .B(AddRoundKeyOutput[61]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n23) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_2_U1 ( .A1(AddRoundKeyOutput[60]), .A2(
        AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U9 ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n23), .A2(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U7 ( .A1(AddRoundKeyOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n23), .A2(
        SubCellInst_LFInst_15_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n20), .A2(
        SubCellInst_LFInst_15_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U4 ( .A1(AddRoundKeyOutput[62]), .A2(
        AddRoundKeyOutput[60]), .ZN(SubCellInst_LFInst_15_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_15_LFInst_3_U3 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U2 ( .A1(AddRoundKeyOutput[60]), .A2(
        AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n26), .A2(
        SubCellInst_LFInst_15_LFInst_3_n25), .ZN(Red_MCInst_MC0_v0_1[0]) );
  BUF_X1 MCInst_MC0_U2 ( .A(ShiftRowsOutput[28]), .Z(MCInst_MC0_v2_3[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U2 ( .A(MCInst_MC0_v0_2Inst_0_n3), .B(
        Red_MCInst_MC0_v0_1[0]), .ZN(MCInst_MC0_v0_2[0]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .ZN(MCInst_MC0_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v1_1Inst_0_U1 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .Z(MCInst_MC0_v1_1[0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U2 ( .A(MCInst_MC0_v1_2Inst_0_n3), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_v1_2[0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v2_1Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(MCInst_MC0_v2_1[0]) );
  XOR2_X1 MCInst_MC0_v2_2Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(MCInst_MC0_v2_2[0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U3 ( .A(MCInst_MC0_v2_3Inst_0_n6), .B(
        MCInst_MC0_v2_3Inst_0_n5), .ZN(MCInst_MC0_v2_3[0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC0_v2_3Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC0_v3_1Inst_0_U1 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_v3_1[0]) );
  XOR2_X1 MCInst_MC0_v3_2Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_v3_2[0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U2 ( .A(MCInst_MC0_v3_3Inst_0_n3), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(MCInst_MC0_v3_3[0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(MCInst_MC0_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v0_0Inst_1_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_0[1]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_1_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v0_3[3]), .Z(MCInst_MC0_v0_1[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U2 ( .A(MCInst_MC0_v0_2Inst_1_n3), .B(
        Red_MCInst_MC0_v0_1[0]), .ZN(MCInst_MC0_v0_2[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .ZN(MCInst_MC0_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_3[1]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[3]), .Z(MCInst_MC0_v1_1[1]) );
  XOR2_X1 MCInst_MC0_v1_2Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .Z(MCInst_MC0_v1_2[1]) );
  XOR2_X1 MCInst_MC0_v1_3Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_1[2]), .Z(MCInst_MC0_v1_3[1]) );
  XOR2_X1 MCInst_MC0_v2_0Inst_1_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(MCInst_MC0_v2_0[1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U2 ( .A(MCInst_MC0_v2_1Inst_1_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_1[1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U3 ( .A(MCInst_MC0_v2_2Inst_1_n6), .B(
        MCInst_MC0_v2_2Inst_1_n5), .ZN(MCInst_MC0_v2_2[1]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC0_v2_2Inst_1_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC0_v3_0Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_v3_0[1]) );
  XOR2_X1 MCInst_MC0_v3_1Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_v3_1[1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U2 ( .A(MCInst_MC0_v3_3Inst_1_n3), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(MCInst_MC0_v3_3[1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .ZN(MCInst_MC0_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_0[2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_2_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_1[2]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_2[2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U2 ( .A(MCInst_MC0_v1_1Inst_2_n3), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_v1_1[2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U2 ( .A(MCInst_MC0_v1_2Inst_2_n3), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_v1_2[2]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U2 ( .A(MCInst_MC0_v2_1Inst_2_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_1[2]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U2 ( .A(MCInst_MC0_v2_2Inst_2_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_2[2]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC0_v2_3Inst_2_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_3[2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U2 ( .A(MCInst_MC0_v3_1Inst_2_n3), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(MCInst_MC0_v3_1[2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(MCInst_MC0_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC0_v3_3Inst_2_U1 ( .A(Red_MCInst_MC0_v3_3[2]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_v3_3[2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_3_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_1[3]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_3_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .Z(MCInst_MC0_v0_2[3]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_3_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        MCInst_MC0_v1_3[3]), .Z(MCInst_MC0_v1_1[3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U3 ( .A(MCInst_MC0_v1_2Inst_3_n6), .B(
        MCInst_MC0_v1_2Inst_3_n5), .ZN(MCInst_MC0_v1_2[3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U2 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC0_v1_2Inst_3_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .Z(MCInst_MC0_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC0_v2_1Inst_3_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(MCInst_MC0_v2_1[3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U2 ( .A(MCInst_MC0_v2_2Inst_3_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_2[3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U2 ( .A(MCInst_MC0_v2_3Inst_3_n3), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_3[3]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .ZN(MCInst_MC0_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC0_v3_1Inst_3_U1 ( .A(Red_MCInst_MC0_v3_3[2]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_v3_1[3]) );
  XOR2_X1 MCInst_MC0_v3_3Inst_3_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_v3_3[3]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_0_n8), .B(MCInst_MC0_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[60]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_2[1]), .B(
        MCInst_MC0_v1_0_0_), .ZN(MCInst_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_1_n8), .B(MCInst_MC0_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[61]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_0[1]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_0[1]), .B(
        MCInst_MC0_v3_0[1]), .Z(MCInst_MC0_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_2_n8), .B(MCInst_MC0_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[62]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_0[2]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_3_n8), .B(MCInst_MC0_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[63]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_0_n8), .B(MCInst_MC0_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[44]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_1[0]), .B(
        MCInst_MC0_v1_1[0]), .ZN(MCInst_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_1[0]), .Z(MCInst_MC0_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_1_n8), .B(MCInst_MC0_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[45]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v1_1[1]), .ZN(MCInst_MC0_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_1[1]), .B(
        MCInst_MC0_v3_1[1]), .Z(MCInst_MC0_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_2_n8), .B(MCInst_MC0_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[46]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_1[2]), .B(
        MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_1[2]), .B(
        MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_3_n8), .B(MCInst_MC0_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[47]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_1[3]), .B(
        MCInst_MC0_v1_1[3]), .ZN(MCInst_MC0_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_1[3]), .B(
        MCInst_MC0_v3_1[3]), .Z(MCInst_MC0_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_0_n8), .B(MCInst_MC0_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[28]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_2[0]), .B(
        MCInst_MC0_v1_2[0]), .ZN(MCInst_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_2[0]), .B(
        MCInst_MC0_v3_2[0]), .Z(MCInst_MC0_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_1_n8), .B(MCInst_MC0_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[29]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_2[1]), .B(
        MCInst_MC0_v1_2[1]), .ZN(MCInst_MC0_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_2[1]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_2_n8), .B(MCInst_MC0_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[30]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_2[2]), .B(
        MCInst_MC0_v1_2[2]), .ZN(MCInst_MC0_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_2[2]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_3_n8), .B(MCInst_MC0_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[31]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_2[3]), .B(
        MCInst_MC0_v1_2[3]), .ZN(MCInst_MC0_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_2[3]), .B(
        MCInst_MC0_v3_2[3]), .Z(MCInst_MC0_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_0_n8), .B(MCInst_MC0_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[12]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_3[0]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_1[0]), .B(
        MCInst_MC0_v3_3[0]), .Z(MCInst_MC0_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_1_n8), .B(MCInst_MC0_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[13]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v1_3[1]), .ZN(MCInst_MC0_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_3[1]), .B(
        MCInst_MC0_v3_3[1]), .Z(MCInst_MC0_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_2_n8), .B(MCInst_MC0_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[14]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_3[2]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_3_n8), .B(MCInst_MC0_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[15]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_3[3]), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v3_3[3]), .Z(MCInst_MC0_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst_MC1_U2 ( .A(ShiftRowsOutput[24]), .Z(MCInst_MC1_v2_3[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U2 ( .A(MCInst_MC1_v0_2Inst_0_n3), .B(
        Red_MCInst_MC1_v0_1[0]), .ZN(MCInst_MC1_v0_2[0]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .ZN(MCInst_MC1_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v1_1Inst_0_U1 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .Z(MCInst_MC1_v1_1[0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U2 ( .A(MCInst_MC1_v1_2Inst_0_n3), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_v1_2[0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v2_1Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(MCInst_MC1_v2_1[0]) );
  XOR2_X1 MCInst_MC1_v2_2Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(MCInst_MC1_v2_2[0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U3 ( .A(MCInst_MC1_v2_3Inst_0_n6), .B(
        MCInst_MC1_v2_3Inst_0_n5), .ZN(MCInst_MC1_v2_3[0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC1_v2_3Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC1_v3_1Inst_0_U1 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_v3_1[0]) );
  XOR2_X1 MCInst_MC1_v3_2Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_v3_2[0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U2 ( .A(MCInst_MC1_v3_3Inst_0_n3), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(MCInst_MC1_v3_3[0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(MCInst_MC1_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v0_0Inst_1_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_0[1]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_1_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v0_3[3]), .Z(MCInst_MC1_v0_1[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U2 ( .A(MCInst_MC1_v0_2Inst_1_n3), .B(
        Red_MCInst_MC1_v0_1[0]), .ZN(MCInst_MC1_v0_2[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .ZN(MCInst_MC1_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_3[1]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[3]), .Z(MCInst_MC1_v1_1[1]) );
  XOR2_X1 MCInst_MC1_v1_2Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .Z(MCInst_MC1_v1_2[1]) );
  XOR2_X1 MCInst_MC1_v1_3Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_1[2]), .Z(MCInst_MC1_v1_3[1]) );
  XOR2_X1 MCInst_MC1_v2_0Inst_1_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(MCInst_MC1_v2_0[1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U2 ( .A(MCInst_MC1_v2_1Inst_1_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_1[1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U3 ( .A(MCInst_MC1_v2_2Inst_1_n6), .B(
        MCInst_MC1_v2_2Inst_1_n5), .ZN(MCInst_MC1_v2_2[1]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC1_v2_2Inst_1_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC1_v3_0Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_v3_0[1]) );
  XOR2_X1 MCInst_MC1_v3_1Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_v3_1[1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U2 ( .A(MCInst_MC1_v3_3Inst_1_n3), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(MCInst_MC1_v3_3[1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .ZN(MCInst_MC1_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_0[2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_2_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_1[2]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_2[2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U2 ( .A(MCInst_MC1_v1_1Inst_2_n3), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_v1_1[2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U2 ( .A(MCInst_MC1_v1_2Inst_2_n3), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_v1_2[2]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U2 ( .A(MCInst_MC1_v2_1Inst_2_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_1[2]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U2 ( .A(MCInst_MC1_v2_2Inst_2_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_2[2]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC1_v2_3Inst_2_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_3[2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U2 ( .A(MCInst_MC1_v3_1Inst_2_n3), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(MCInst_MC1_v3_1[2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(MCInst_MC1_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC1_v3_3Inst_2_U1 ( .A(Red_MCInst_MC1_v3_3[2]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_v3_3[2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_3_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_1[3]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_3_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .Z(MCInst_MC1_v0_2[3]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_3_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        MCInst_MC1_v1_3[3]), .Z(MCInst_MC1_v1_1[3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U3 ( .A(MCInst_MC1_v1_2Inst_3_n6), .B(
        MCInst_MC1_v1_2Inst_3_n5), .ZN(MCInst_MC1_v1_2[3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U2 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC1_v1_2Inst_3_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .Z(MCInst_MC1_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC1_v2_1Inst_3_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(MCInst_MC1_v2_1[3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U2 ( .A(MCInst_MC1_v2_2Inst_3_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_2[3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U2 ( .A(MCInst_MC1_v2_3Inst_3_n3), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_3[3]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .ZN(MCInst_MC1_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC1_v3_1Inst_3_U1 ( .A(Red_MCInst_MC1_v3_3[2]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_v3_1[3]) );
  XOR2_X1 MCInst_MC1_v3_3Inst_3_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_v3_3[3]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_0_n8), .B(MCInst_MC1_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[56]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_2[1]), .B(
        MCInst_MC1_v1_0_0_), .ZN(MCInst_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_1_n8), .B(MCInst_MC1_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[57]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_0[1]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_0[1]), .B(
        MCInst_MC1_v3_0[1]), .Z(MCInst_MC1_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_2_n8), .B(MCInst_MC1_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[58]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_0[2]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_3_n8), .B(MCInst_MC1_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[59]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_0_n8), .B(MCInst_MC1_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[40]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_1[0]), .B(
        MCInst_MC1_v1_1[0]), .ZN(MCInst_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_1[0]), .Z(MCInst_MC1_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_1_n8), .B(MCInst_MC1_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[41]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v1_1[1]), .ZN(MCInst_MC1_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_1[1]), .B(
        MCInst_MC1_v3_1[1]), .Z(MCInst_MC1_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_2_n8), .B(MCInst_MC1_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[42]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_1[2]), .B(
        MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_1[2]), .B(
        MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_3_n8), .B(MCInst_MC1_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[43]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_1[3]), .B(
        MCInst_MC1_v1_1[3]), .ZN(MCInst_MC1_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_1[3]), .B(
        MCInst_MC1_v3_1[3]), .Z(MCInst_MC1_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_0_n8), .B(MCInst_MC1_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[24]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_2[0]), .B(
        MCInst_MC1_v1_2[0]), .ZN(MCInst_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_2[0]), .B(
        MCInst_MC1_v3_2[0]), .Z(MCInst_MC1_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_1_n8), .B(MCInst_MC1_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[25]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_2[1]), .B(
        MCInst_MC1_v1_2[1]), .ZN(MCInst_MC1_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_2[1]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_2_n8), .B(MCInst_MC1_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[26]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_2[2]), .B(
        MCInst_MC1_v1_2[2]), .ZN(MCInst_MC1_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_2[2]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_3_n8), .B(MCInst_MC1_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[27]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_2[3]), .B(
        MCInst_MC1_v1_2[3]), .ZN(MCInst_MC1_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_2[3]), .B(
        MCInst_MC1_v3_2[3]), .Z(MCInst_MC1_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_0_n8), .B(MCInst_MC1_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[8]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_3[0]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_1[0]), .B(
        MCInst_MC1_v3_3[0]), .Z(MCInst_MC1_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_1_n8), .B(MCInst_MC1_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[9]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v1_3[1]), .ZN(MCInst_MC1_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_3[1]), .B(
        MCInst_MC1_v3_3[1]), .Z(MCInst_MC1_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_2_n8), .B(MCInst_MC1_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[10]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_3[2]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_3_n8), .B(MCInst_MC1_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[11]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_3[3]), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v3_3[3]), .Z(MCInst_MC1_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst_MC2_U2 ( .A(ShiftRowsOutput[20]), .Z(MCInst_MC2_v2_3[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U2 ( .A(MCInst_MC2_v0_2Inst_0_n3), .B(
        Red_MCInst_MC2_v0_1[0]), .ZN(MCInst_MC2_v0_2[0]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .ZN(MCInst_MC2_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v1_1Inst_0_U1 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .Z(MCInst_MC2_v1_1[0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U2 ( .A(MCInst_MC2_v1_2Inst_0_n3), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_v1_2[0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v2_1Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(MCInst_MC2_v2_1[0]) );
  XOR2_X1 MCInst_MC2_v2_2Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(MCInst_MC2_v2_2[0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U3 ( .A(MCInst_MC2_v2_3Inst_0_n6), .B(
        MCInst_MC2_v2_3Inst_0_n5), .ZN(MCInst_MC2_v2_3[0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC2_v2_3Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC2_v3_1Inst_0_U1 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_v3_1[0]) );
  XOR2_X1 MCInst_MC2_v3_2Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_v3_2[0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U2 ( .A(MCInst_MC2_v3_3Inst_0_n3), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(MCInst_MC2_v3_3[0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(MCInst_MC2_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v0_0Inst_1_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_0[1]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_1_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v0_3[3]), .Z(MCInst_MC2_v0_1[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U2 ( .A(MCInst_MC2_v0_2Inst_1_n3), .B(
        Red_MCInst_MC2_v0_1[0]), .ZN(MCInst_MC2_v0_2[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .ZN(MCInst_MC2_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_3[1]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[3]), .Z(MCInst_MC2_v1_1[1]) );
  XOR2_X1 MCInst_MC2_v1_2Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .Z(MCInst_MC2_v1_2[1]) );
  XOR2_X1 MCInst_MC2_v1_3Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_1[2]), .Z(MCInst_MC2_v1_3[1]) );
  XOR2_X1 MCInst_MC2_v2_0Inst_1_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(MCInst_MC2_v2_0[1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U2 ( .A(MCInst_MC2_v2_1Inst_1_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_1[1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U3 ( .A(MCInst_MC2_v2_2Inst_1_n6), .B(
        MCInst_MC2_v2_2Inst_1_n5), .ZN(MCInst_MC2_v2_2[1]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC2_v2_2Inst_1_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC2_v3_0Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_v3_0[1]) );
  XOR2_X1 MCInst_MC2_v3_1Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_v3_1[1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U2 ( .A(MCInst_MC2_v3_3Inst_1_n3), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(MCInst_MC2_v3_3[1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .ZN(MCInst_MC2_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_0[2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_2_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_1[2]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_2[2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U2 ( .A(MCInst_MC2_v1_1Inst_2_n3), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_v1_1[2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U2 ( .A(MCInst_MC2_v1_2Inst_2_n3), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_v1_2[2]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U2 ( .A(MCInst_MC2_v2_1Inst_2_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_1[2]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U2 ( .A(MCInst_MC2_v2_2Inst_2_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_2[2]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC2_v2_3Inst_2_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_3[2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U2 ( .A(MCInst_MC2_v3_1Inst_2_n3), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(MCInst_MC2_v3_1[2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(MCInst_MC2_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC2_v3_3Inst_2_U1 ( .A(Red_MCInst_MC2_v3_3[2]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_v3_3[2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_3_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_1[3]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_3_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .Z(MCInst_MC2_v0_2[3]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_3_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        MCInst_MC2_v1_3[3]), .Z(MCInst_MC2_v1_1[3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U3 ( .A(MCInst_MC2_v1_2Inst_3_n6), .B(
        MCInst_MC2_v1_2Inst_3_n5), .ZN(MCInst_MC2_v1_2[3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U2 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC2_v1_2Inst_3_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .Z(MCInst_MC2_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC2_v2_1Inst_3_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(MCInst_MC2_v2_1[3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U2 ( .A(MCInst_MC2_v2_2Inst_3_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_2[3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U2 ( .A(MCInst_MC2_v2_3Inst_3_n3), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_3[3]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .ZN(MCInst_MC2_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC2_v3_1Inst_3_U1 ( .A(Red_MCInst_MC2_v3_3[2]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_v3_1[3]) );
  XOR2_X1 MCInst_MC2_v3_3Inst_3_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_v3_3[3]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_0_n8), .B(MCInst_MC2_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[52]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_2[1]), .B(
        MCInst_MC2_v1_0_0_), .ZN(MCInst_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_1_n8), .B(MCInst_MC2_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[53]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_0[1]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_0[1]), .B(
        MCInst_MC2_v3_0[1]), .Z(MCInst_MC2_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_2_n8), .B(MCInst_MC2_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[54]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_0[2]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_3_n8), .B(MCInst_MC2_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[55]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_0_n8), .B(MCInst_MC2_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[36]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_1[0]), .B(
        MCInst_MC2_v1_1[0]), .ZN(MCInst_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_1[0]), .Z(MCInst_MC2_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_1_n8), .B(MCInst_MC2_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[37]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v1_1[1]), .ZN(MCInst_MC2_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_1[1]), .B(
        MCInst_MC2_v3_1[1]), .Z(MCInst_MC2_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_2_n8), .B(MCInst_MC2_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[38]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_1[2]), .B(
        MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_1[2]), .B(
        MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_3_n8), .B(MCInst_MC2_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[39]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_1[3]), .B(
        MCInst_MC2_v1_1[3]), .ZN(MCInst_MC2_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_1[3]), .B(
        MCInst_MC2_v3_1[3]), .Z(MCInst_MC2_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_0_n8), .B(MCInst_MC2_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[20]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_2[0]), .B(
        MCInst_MC2_v1_2[0]), .ZN(MCInst_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_2[0]), .B(
        MCInst_MC2_v3_2[0]), .Z(MCInst_MC2_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_1_n8), .B(MCInst_MC2_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[21]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_2[1]), .B(
        MCInst_MC2_v1_2[1]), .ZN(MCInst_MC2_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_2[1]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_2_n8), .B(MCInst_MC2_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[22]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_2[2]), .B(
        MCInst_MC2_v1_2[2]), .ZN(MCInst_MC2_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_2[2]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_3_n8), .B(MCInst_MC2_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[23]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_2[3]), .B(
        MCInst_MC2_v1_2[3]), .ZN(MCInst_MC2_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_2[3]), .B(
        MCInst_MC2_v3_2[3]), .Z(MCInst_MC2_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_0_n8), .B(MCInst_MC2_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[4]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_3[0]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_1[0]), .B(
        MCInst_MC2_v3_3[0]), .Z(MCInst_MC2_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_1_n8), .B(MCInst_MC2_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[5]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v1_3[1]), .ZN(MCInst_MC2_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_3[1]), .B(
        MCInst_MC2_v3_3[1]), .Z(MCInst_MC2_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_2_n8), .B(MCInst_MC2_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[6]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_3[2]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_3_n8), .B(MCInst_MC2_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[7]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_3[3]), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v3_3[3]), .Z(MCInst_MC2_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst_MC3_U2 ( .A(ShiftRowsOutput[16]), .Z(MCInst_MC3_v2_3[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U2 ( .A(MCInst_MC3_v0_2Inst_0_n3), .B(
        Red_MCInst_MC3_v0_1[0]), .ZN(MCInst_MC3_v0_2[0]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .ZN(MCInst_MC3_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v1_1Inst_0_U1 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .Z(MCInst_MC3_v1_1[0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U2 ( .A(MCInst_MC3_v1_2Inst_0_n3), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_v1_2[0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v2_1Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(MCInst_MC3_v2_1[0]) );
  XOR2_X1 MCInst_MC3_v2_2Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(MCInst_MC3_v2_2[0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U3 ( .A(MCInst_MC3_v2_3Inst_0_n6), .B(
        MCInst_MC3_v2_3Inst_0_n5), .ZN(MCInst_MC3_v2_3[0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC3_v2_3Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC3_v3_1Inst_0_U1 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_v3_1[0]) );
  XOR2_X1 MCInst_MC3_v3_2Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_v3_2[0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U2 ( .A(MCInst_MC3_v3_3Inst_0_n3), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(MCInst_MC3_v3_3[0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(MCInst_MC3_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v0_0Inst_1_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_0[1]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_1_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v0_3[3]), .Z(MCInst_MC3_v0_1[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U2 ( .A(MCInst_MC3_v0_2Inst_1_n3), .B(
        Red_MCInst_MC3_v0_1[0]), .ZN(MCInst_MC3_v0_2[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .ZN(MCInst_MC3_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_3[1]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[3]), .Z(MCInst_MC3_v1_1[1]) );
  XOR2_X1 MCInst_MC3_v1_2Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .Z(MCInst_MC3_v1_2[1]) );
  XOR2_X1 MCInst_MC3_v1_3Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_1[2]), .Z(MCInst_MC3_v1_3[1]) );
  XOR2_X1 MCInst_MC3_v2_0Inst_1_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(MCInst_MC3_v2_0[1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U2 ( .A(MCInst_MC3_v2_1Inst_1_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_1[1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U3 ( .A(MCInst_MC3_v2_2Inst_1_n6), .B(
        MCInst_MC3_v2_2Inst_1_n5), .ZN(MCInst_MC3_v2_2[1]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC3_v2_2Inst_1_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC3_v3_0Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_v3_0[1]) );
  XOR2_X1 MCInst_MC3_v3_1Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_v3_1[1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U2 ( .A(MCInst_MC3_v3_3Inst_1_n3), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(MCInst_MC3_v3_3[1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .ZN(MCInst_MC3_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_0[2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_2_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_1[2]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_2[2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U2 ( .A(MCInst_MC3_v1_1Inst_2_n3), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_v1_1[2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U2 ( .A(MCInst_MC3_v1_2Inst_2_n3), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_v1_2[2]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U2 ( .A(MCInst_MC3_v2_1Inst_2_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_1[2]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U2 ( .A(MCInst_MC3_v2_2Inst_2_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_2[2]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC3_v2_3Inst_2_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_3[2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U2 ( .A(MCInst_MC3_v3_1Inst_2_n3), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(MCInst_MC3_v3_1[2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(MCInst_MC3_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC3_v3_3Inst_2_U1 ( .A(Red_MCInst_MC3_v3_3[2]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_v3_3[2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_3_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_1[3]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_3_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .Z(MCInst_MC3_v0_2[3]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_3_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        MCInst_MC3_v1_3[3]), .Z(MCInst_MC3_v1_1[3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U3 ( .A(MCInst_MC3_v1_2Inst_3_n6), .B(
        MCInst_MC3_v1_2Inst_3_n5), .ZN(MCInst_MC3_v1_2[3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U2 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC3_v1_2Inst_3_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .Z(MCInst_MC3_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC3_v2_1Inst_3_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(MCInst_MC3_v2_1[3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U2 ( .A(MCInst_MC3_v2_2Inst_3_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_2[3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U2 ( .A(MCInst_MC3_v2_3Inst_3_n3), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_3[3]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .ZN(MCInst_MC3_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC3_v3_1Inst_3_U1 ( .A(Red_MCInst_MC3_v3_3[2]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_v3_1[3]) );
  XOR2_X1 MCInst_MC3_v3_3Inst_3_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_v3_3[3]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_0_n8), .B(MCInst_MC3_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[48]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_2[1]), .B(
        MCInst_MC3_v1_0_0_), .ZN(MCInst_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_1_n8), .B(MCInst_MC3_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[49]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_0[1]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_0[1]), .B(
        MCInst_MC3_v3_0[1]), .Z(MCInst_MC3_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_2_n8), .B(MCInst_MC3_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[50]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_0[2]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_3_n8), .B(MCInst_MC3_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[51]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_0_n8), .B(MCInst_MC3_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[32]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_1[0]), .B(
        MCInst_MC3_v1_1[0]), .ZN(MCInst_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_1[0]), .Z(MCInst_MC3_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_1_n8), .B(MCInst_MC3_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[33]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v1_1[1]), .ZN(MCInst_MC3_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_1[1]), .B(
        MCInst_MC3_v3_1[1]), .Z(MCInst_MC3_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_2_n8), .B(MCInst_MC3_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[34]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_1[2]), .B(
        MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_1[2]), .B(
        MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_3_n8), .B(MCInst_MC3_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[35]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_1[3]), .B(
        MCInst_MC3_v1_1[3]), .ZN(MCInst_MC3_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_1[3]), .B(
        MCInst_MC3_v3_1[3]), .Z(MCInst_MC3_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_0_n8), .B(MCInst_MC3_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[16]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_2[0]), .B(
        MCInst_MC3_v1_2[0]), .ZN(MCInst_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_2[0]), .B(
        MCInst_MC3_v3_2[0]), .Z(MCInst_MC3_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_1_n8), .B(MCInst_MC3_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[17]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_2[1]), .B(
        MCInst_MC3_v1_2[1]), .ZN(MCInst_MC3_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_2[1]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_2_n8), .B(MCInst_MC3_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[18]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_2[2]), .B(
        MCInst_MC3_v1_2[2]), .ZN(MCInst_MC3_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_2[2]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_3_n8), .B(MCInst_MC3_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[19]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_2[3]), .B(
        MCInst_MC3_v1_2[3]), .ZN(MCInst_MC3_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_2[3]), .B(
        MCInst_MC3_v3_2[3]), .Z(MCInst_MC3_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_0_n8), .B(MCInst_MC3_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[0]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_3[0]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_1[0]), .B(
        MCInst_MC3_v3_3[0]), .Z(MCInst_MC3_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_1_n8), .B(MCInst_MC3_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[1]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v1_3[1]), .ZN(MCInst_MC3_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_3[1]), .B(
        MCInst_MC3_v3_3[1]), .Z(MCInst_MC3_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_2_n8), .B(MCInst_MC3_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[2]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_3[2]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_3_n8), .B(MCInst_MC3_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[3]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_3[3]), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v3_3[3]), .Z(MCInst_MC3_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n3), .B(Plaintext[2]), .ZN(
        Red_Plaintext[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Plaintext[0]), .B(
        Plaintext[1]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_1_n3), .B(Plaintext[3]), .ZN(
        Red_Plaintext[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U1 ( .A(Plaintext[0]), .B(
        Plaintext[1]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_2_n3), .B(Plaintext[3]), .ZN(
        Red_Plaintext[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U1 ( .A(Plaintext[1]), .B(
        Plaintext[2]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n3), .B(Plaintext[6]), .ZN(
        Red_Plaintext[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Plaintext[4]), .B(
        Plaintext[5]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_1_n3), .B(Plaintext[7]), .ZN(
        Red_Plaintext[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U1 ( .A(Plaintext[4]), .B(
        Plaintext[5]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_2_n3), .B(Plaintext[7]), .ZN(
        Red_Plaintext[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U1 ( .A(Plaintext[5]), .B(
        Plaintext[6]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n3), .B(Plaintext[10]), .ZN(
        Red_Plaintext[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Plaintext[8]), .B(
        Plaintext[9]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_1_n3), .B(Plaintext[11]), .ZN(
        Red_Plaintext[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U1 ( .A(Plaintext[8]), .B(
        Plaintext[9]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_2_n3), .B(Plaintext[11]), .ZN(
        Red_Plaintext[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U1 ( .A(Plaintext[9]), .B(
        Plaintext[10]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n3), .B(Plaintext[14]), .ZN(
        Red_Plaintext[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Plaintext[12]), .B(
        Plaintext[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_1_n3), .B(Plaintext[15]), .ZN(
        Red_Plaintext[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U1 ( .A(Plaintext[12]), .B(
        Plaintext[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_2_n3), .B(Plaintext[15]), .ZN(
        Red_Plaintext[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U1 ( .A(Plaintext[13]), .B(
        Plaintext[14]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n3), .B(Plaintext[18]), .ZN(
        Red_Plaintext[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Plaintext[16]), .B(
        Plaintext[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_1_n3), .B(Plaintext[19]), .ZN(
        Red_Plaintext[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U1 ( .A(Plaintext[16]), .B(
        Plaintext[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_2_n3), .B(Plaintext[19]), .ZN(
        Red_Plaintext[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U1 ( .A(Plaintext[17]), .B(
        Plaintext[18]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n3), .B(Plaintext[22]), .ZN(
        Red_Plaintext[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Plaintext[20]), .B(
        Plaintext[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_1_n3), .B(Plaintext[23]), .ZN(
        Red_Plaintext[16]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U1 ( .A(Plaintext[20]), .B(
        Plaintext[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_2_n3), .B(Plaintext[23]), .ZN(
        Red_Plaintext[17]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U1 ( .A(Plaintext[21]), .B(
        Plaintext[22]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n3), .B(Plaintext[26]), .ZN(
        Red_Plaintext[18]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Plaintext[24]), .B(
        Plaintext[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_1_n3), .B(Plaintext[27]), .ZN(
        Red_Plaintext[19]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U1 ( .A(Plaintext[24]), .B(
        Plaintext[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_2_n3), .B(Plaintext[27]), .ZN(
        Red_Plaintext[20]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U1 ( .A(Plaintext[25]), .B(
        Plaintext[26]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n3), .B(Plaintext[30]), .ZN(
        Red_Plaintext[21]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Plaintext[28]), .B(
        Plaintext[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_1_n3), .B(Plaintext[31]), .ZN(
        Red_Plaintext[22]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U1 ( .A(Plaintext[28]), .B(
        Plaintext[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_2_n3), .B(Plaintext[31]), .ZN(
        Red_Plaintext[23]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U1 ( .A(Plaintext[29]), .B(
        Plaintext[30]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n3), .B(Plaintext[34]), .ZN(
        Red_Plaintext[24]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Plaintext[32]), .B(
        Plaintext[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_1_n3), .B(Plaintext[35]), .ZN(
        Red_Plaintext[25]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U1 ( .A(Plaintext[32]), .B(
        Plaintext[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_2_n3), .B(Plaintext[35]), .ZN(
        Red_Plaintext[26]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U1 ( .A(Plaintext[33]), .B(
        Plaintext[34]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n3), .B(Plaintext[38]), .ZN(
        Red_Plaintext[27]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Plaintext[36]), .B(
        Plaintext[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_1_n3), .B(Plaintext[39]), .ZN(
        Red_Plaintext[28]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U1 ( .A(Plaintext[36]), .B(
        Plaintext[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_2_n3), .B(Plaintext[39]), .ZN(
        Red_Plaintext[29]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U1 ( .A(Plaintext[37]), .B(
        Plaintext[38]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n3), .B(Plaintext[42]), .ZN(
        Red_Plaintext[30]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Plaintext[40]), .B(
        Plaintext[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_1_n3), .B(Plaintext[43]), .ZN(
        Red_Plaintext[31]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U1 ( .A(Plaintext[40]), .B(
        Plaintext[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_2_n3), .B(Plaintext[43]), .ZN(
        Red_Plaintext[32]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U1 ( .A(Plaintext[41]), .B(
        Plaintext[42]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n3), .B(Plaintext[46]), .ZN(
        Red_Plaintext[33]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Plaintext[44]), .B(
        Plaintext[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_1_n3), .B(Plaintext[47]), .ZN(
        Red_Plaintext[34]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U1 ( .A(Plaintext[44]), .B(
        Plaintext[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_2_n3), .B(Plaintext[47]), .ZN(
        Red_Plaintext[35]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U1 ( .A(Plaintext[45]), .B(
        Plaintext[46]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n3), .B(Plaintext[50]), .ZN(
        Red_Plaintext[36]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Plaintext[48]), .B(
        Plaintext[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_1_n3), .B(Plaintext[51]), .ZN(
        Red_Plaintext[37]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U1 ( .A(Plaintext[48]), .B(
        Plaintext[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_2_n3), .B(Plaintext[51]), .ZN(
        Red_Plaintext[38]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U1 ( .A(Plaintext[49]), .B(
        Plaintext[50]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n3), .B(Plaintext[54]), .ZN(
        Red_Plaintext[39]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Plaintext[52]), .B(
        Plaintext[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_1_n3), .B(Plaintext[55]), .ZN(
        Red_Plaintext[40]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U1 ( .A(Plaintext[52]), .B(
        Plaintext[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_2_n3), .B(Plaintext[55]), .ZN(
        Red_Plaintext[41]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U1 ( .A(Plaintext[53]), .B(
        Plaintext[54]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n3), .B(Plaintext[58]), .ZN(
        Red_Plaintext[42]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Plaintext[56]), .B(
        Plaintext[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_1_n3), .B(Plaintext[59]), .ZN(
        Red_Plaintext[43]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U1 ( .A(Plaintext[56]), .B(
        Plaintext[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_2_n3), .B(Plaintext[59]), .ZN(
        Red_Plaintext[44]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U1 ( .A(Plaintext[57]), .B(
        Plaintext[58]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n3), .B(Plaintext[62]), .ZN(
        Red_Plaintext[45]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Plaintext[60]), .B(
        Plaintext[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_1_n3), .B(Plaintext[63]), .ZN(
        Red_Plaintext[46]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U1 ( .A(Plaintext[60]), .B(
        Plaintext[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_2_n3), .B(Plaintext[63]), .ZN(
        Red_Plaintext[47]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U1 ( .A(Plaintext[61]), .B(
        Plaintext[62]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_2_n3) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_0_U1 ( .A(Red_Plaintext[0]), .B(
        Red_RoundKey[0]), .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_1_U1 ( .A(Red_Plaintext[1]), .B(
        Red_RoundKey[1]), .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_2_U1 ( .A(Red_Plaintext[2]), .B(
        Red_RoundKey[2]), .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_0_U1 ( .A(Red_Plaintext[3]), .B(
        Red_RoundKey[3]), .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_1_U1 ( .A(Red_Plaintext[4]), .B(
        Red_RoundKey[4]), .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_2_U1 ( .A(Red_Plaintext[5]), .B(
        Red_RoundKey[5]), .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_0_U1 ( .A(Red_Plaintext[6]), .B(
        Red_RoundKey[6]), .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_1_U1 ( .A(Red_Plaintext[7]), .B(
        Red_RoundKey[7]), .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_2_U1 ( .A(Red_Plaintext[8]), .B(
        Red_RoundKey[8]), .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_0_U1 ( .A(Red_Plaintext[9]), .B(
        Red_RoundKey[9]), .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_1_U1 ( .A(Red_Plaintext[10]), .B(
        Red_RoundKey[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_2_U1 ( .A(Red_Plaintext[11]), .B(
        Red_RoundKey[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_0_U1 ( .A(Red_Plaintext[12]), .B(
        Red_RoundKey[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_1_U1 ( .A(Red_Plaintext[13]), .B(
        Red_RoundKey[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_2_U1 ( .A(Red_Plaintext[14]), .B(
        Red_RoundKey[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_0_U1 ( .A(Red_Plaintext[15]), .B(
        Red_RoundKey[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_1_U1 ( .A(Red_Plaintext[16]), .B(
        Red_RoundKey[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_2_U1 ( .A(Red_Plaintext[17]), .B(
        Red_RoundKey[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_0_U1 ( .A(Red_Plaintext[18]), .B(
        Red_RoundKey[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_1_U1 ( .A(Red_Plaintext[19]), .B(
        Red_RoundKey[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_2_U1 ( .A(Red_Plaintext[20]), .B(
        Red_RoundKey[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_0_U1 ( .A(Red_Plaintext[21]), .B(
        Red_RoundKey[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_1_U1 ( .A(Red_Plaintext[22]), .B(
        Red_RoundKey[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_2_U1 ( .A(Red_Plaintext[23]), .B(
        Red_RoundKey[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_0_U1 ( .A(Red_Plaintext[24]), .B(
        Red_RoundKey[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_1_U1 ( .A(Red_Plaintext[25]), .B(
        Red_RoundKey[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_2_U1 ( .A(Red_Plaintext[26]), .B(
        Red_RoundKey[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_0_U1 ( .A(Red_Plaintext[27]), .B(
        Red_RoundKey[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_1_U1 ( .A(Red_Plaintext[28]), .B(
        Red_RoundKey[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_2_U1 ( .A(Red_Plaintext[29]), .B(
        Red_RoundKey[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_0_U1 ( .A(Red_Plaintext[30]), .B(
        Red_RoundKey[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_1_U1 ( .A(Red_Plaintext[31]), .B(
        Red_RoundKey[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_2_U1 ( .A(Red_Plaintext[32]), .B(
        Red_RoundKey[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_0_U1 ( .A(Red_Plaintext[33]), .B(
        Red_RoundKey[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_1_U1 ( .A(Red_Plaintext[34]), .B(
        Red_RoundKey[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_2_U1 ( .A(Red_Plaintext[35]), .B(
        Red_RoundKey[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_0_U1 ( .A(Red_Plaintext[36]), .B(
        Red_RoundKey[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_1_U1 ( .A(Red_Plaintext[37]), .B(
        Red_RoundKey[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_2_U1 ( .A(Red_Plaintext[38]), .B(
        Red_RoundKey[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_0_U1 ( .A(Red_Plaintext[39]), .B(
        Red_RoundKey[39]), .Z(Red_AddRoundKeyOutput[39]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_1_U1 ( .A(Red_Plaintext[40]), .B(
        Red_RoundKey[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_2_U1 ( .A(Red_Plaintext[41]), .B(
        Red_RoundKey[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_0_U1 ( .A(Red_Plaintext[42]), .B(
        Red_RoundKey[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_1_U1 ( .A(Red_Plaintext[43]), .B(
        Red_RoundKey[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_2_U1 ( .A(Red_Plaintext[44]), .B(
        Red_RoundKey[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_0_U1 ( .A(Red_Plaintext[45]), .B(
        Red_RoundKey[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_1_U1 ( .A(Red_Plaintext[46]), .B(
        Red_RoundKey[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_2_U1 ( .A(Red_Plaintext[47]), .B(
        Red_RoundKey[47]), .Z(Red_AddRoundKeyOutput[47]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[9]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U4 ( .A1(AddRoundKeyOutput[2]), 
        .A2(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U3 ( .A1(AddRoundKeyOutput[0]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U2 ( .A1(AddRoundKeyOutput[2]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput[1]), 
        .B(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_0_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[10]) );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U2 ( .A1(AddRoundKeyOutput[3]), 
        .A2(AddRoundKeyOutput[2]), .ZN(Red_SubCellInst_LFInst_0_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U1 ( .A1(AddRoundKeyOutput[1]), 
        .A2(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U7 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n17), .A2(
        Red_SubCellInst_LFInst_0_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[11])
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n15), .A2(AddRoundKeyOutput[3]), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n14), .A2(AddRoundKeyOutput[2]), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U4 ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n13), .A2(
        Red_SubCellInst_LFInst_0_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n17) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_2_U2 ( .A(AddRoundKeyOutput[1]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[2]), .Z(Red_SubCellInst_LFInst_0_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[0]) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U4 ( .A1(AddRoundKeyOutput[6]), 
        .A2(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U3 ( .A1(AddRoundKeyOutput[4]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U2 ( .A1(AddRoundKeyOutput[6]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput[5]), 
        .B(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_1_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[1]) );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U2 ( .A1(AddRoundKeyOutput[7]), 
        .A2(AddRoundKeyOutput[6]), .ZN(Red_SubCellInst_LFInst_1_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U1 ( .A1(AddRoundKeyOutput[5]), 
        .A2(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_1_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[2]) );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(AddRoundKeyOutput[5]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U4 ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[4]), .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n13), .A2(AddRoundKeyOutput[7]), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n12), .A2(AddRoundKeyOutput[6]), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U1 ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[3]) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U4 ( .A1(AddRoundKeyOutput[10]), 
        .A2(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U3 ( .A1(AddRoundKeyOutput[8]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U2 ( .A1(AddRoundKeyOutput[10]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput[9]), 
        .B(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_2_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[4]) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U2 ( .A1(AddRoundKeyOutput[11]), 
        .A2(AddRoundKeyOutput[10]), .ZN(Red_SubCellInst_LFInst_2_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U1 ( .A1(AddRoundKeyOutput[9]), 
        .A2(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_2_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[5]) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(AddRoundKeyOutput[9]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U4 ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[8]), .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n13), .A2(AddRoundKeyOutput[11]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n12), .A2(AddRoundKeyOutput[10]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U1 ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[6]) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U4 ( .A1(AddRoundKeyOutput[14]), 
        .A2(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U3 ( .A1(AddRoundKeyOutput[12]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U2 ( .A1(AddRoundKeyOutput[14]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput[13]), 
        .B(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_3_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[7]) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U2 ( .A1(AddRoundKeyOutput[15]), 
        .A2(AddRoundKeyOutput[14]), .ZN(Red_SubCellInst_LFInst_3_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U1 ( .A1(AddRoundKeyOutput[13]), 
        .A2(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_3_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[8]) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(AddRoundKeyOutput[13]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U4 ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[12]), .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n13), .A2(AddRoundKeyOutput[15]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n12), .A2(AddRoundKeyOutput[14]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U1 ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_4_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[18])
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U4 ( .A1(AddRoundKeyOutput[18]), 
        .A2(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(AddRoundKeyOutput[16]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U2 ( .A1(AddRoundKeyOutput[18]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[17]), 
        .B(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_4_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[19]) );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U2 ( .A1(AddRoundKeyOutput[19]), 
        .A2(AddRoundKeyOutput[18]), .ZN(Red_SubCellInst_LFInst_4_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(AddRoundKeyOutput[17]), 
        .A2(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_4_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[20])
         );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U5 ( .A1(AddRoundKeyOutput[17]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U4 ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[16]), .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n13), .A2(AddRoundKeyOutput[19]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n12), .A2(AddRoundKeyOutput[18]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U1 ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_5_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[21])
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U4 ( .A1(AddRoundKeyOutput[22]), 
        .A2(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(AddRoundKeyOutput[20]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U2 ( .A1(AddRoundKeyOutput[22]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[21]), 
        .B(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_5_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[22]) );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U2 ( .A1(AddRoundKeyOutput[23]), 
        .A2(AddRoundKeyOutput[22]), .ZN(Red_SubCellInst_LFInst_5_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(AddRoundKeyOutput[21]), 
        .A2(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_5_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[23])
         );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U5 ( .A1(AddRoundKeyOutput[21]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U4 ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[20]), .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n13), .A2(AddRoundKeyOutput[23]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n12), .A2(AddRoundKeyOutput[22]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U1 ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_6_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[12])
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U4 ( .A1(AddRoundKeyOutput[26]), 
        .A2(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(AddRoundKeyOutput[24]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U2 ( .A1(AddRoundKeyOutput[26]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[25]), 
        .B(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_6_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[13]) );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U2 ( .A1(AddRoundKeyOutput[27]), 
        .A2(AddRoundKeyOutput[26]), .ZN(Red_SubCellInst_LFInst_6_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(AddRoundKeyOutput[25]), 
        .A2(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_6_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[14])
         );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U5 ( .A1(AddRoundKeyOutput[25]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U4 ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[24]), .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n13), .A2(AddRoundKeyOutput[27]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n12), .A2(AddRoundKeyOutput[26]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U1 ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_7_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[15])
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U4 ( .A1(AddRoundKeyOutput[30]), 
        .A2(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(AddRoundKeyOutput[28]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U2 ( .A1(AddRoundKeyOutput[30]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[29]), 
        .B(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_7_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[16]) );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U2 ( .A1(AddRoundKeyOutput[31]), 
        .A2(AddRoundKeyOutput[30]), .ZN(Red_SubCellInst_LFInst_7_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(AddRoundKeyOutput[29]), 
        .A2(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U7 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n17), .A2(
        Red_SubCellInst_LFInst_7_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[17])
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n15), .A2(AddRoundKeyOutput[31]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n14), .A2(AddRoundKeyOutput[30]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U4 ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n13), .A2(
        Red_SubCellInst_LFInst_7_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_2_n17) );
  INV_X1 Red_SubCellInst_LFInst_7_LFInst_2_U2 ( .A(AddRoundKeyOutput[29]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[30]), .Z(Red_SubCellInst_LFInst_7_LFInst_2_n13)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[27])
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U4 ( .A1(AddRoundKeyOutput[34]), 
        .A2(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U3 ( .A1(AddRoundKeyOutput[32]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U2 ( .A1(AddRoundKeyOutput[34]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput[33]), 
        .B(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_8_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[28]) );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(AddRoundKeyOutput[35]), 
        .A2(AddRoundKeyOutput[34]), .ZN(Red_SubCellInst_LFInst_8_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U1 ( .A1(AddRoundKeyOutput[33]), 
        .A2(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_8_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[29])
         );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U5 ( .A1(AddRoundKeyOutput[33]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U4 ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[32]), .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n13), .A2(AddRoundKeyOutput[35]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n12), .A2(AddRoundKeyOutput[34]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U1 ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[30])
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U4 ( .A1(AddRoundKeyOutput[38]), 
        .A2(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U3 ( .A1(AddRoundKeyOutput[36]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U2 ( .A1(AddRoundKeyOutput[38]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput[37]), 
        .B(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_9_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[31]) );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(AddRoundKeyOutput[39]), 
        .A2(AddRoundKeyOutput[38]), .ZN(Red_SubCellInst_LFInst_9_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U1 ( .A1(AddRoundKeyOutput[37]), 
        .A2(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n11), .A2(
        Red_SubCellInst_LFInst_9_LFInst_2_n13), .ZN(Red_ShiftRowsOutput[32])
         );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(AddRoundKeyOutput[37]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_2_n13) );
  XNOR2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U4 ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[36]), .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n10), .A2(AddRoundKeyOutput[39]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n11) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n9), .A2(AddRoundKeyOutput[38]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n10) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U1 ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[33])
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U4 ( .A1(AddRoundKeyOutput[42]), 
        .A2(AddRoundKeyOutput[43]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U3 ( .A1(AddRoundKeyOutput[40]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U2 ( .A1(AddRoundKeyOutput[42]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput[41]), 
        .B(AddRoundKeyOutput[43]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_10_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[34])
         );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(AddRoundKeyOutput[43]), 
        .A2(AddRoundKeyOutput[42]), .ZN(Red_SubCellInst_LFInst_10_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U1 ( .A1(AddRoundKeyOutput[41]), 
        .A2(AddRoundKeyOutput[43]), .ZN(Red_SubCellInst_LFInst_10_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_10_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[35])
         );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(AddRoundKeyOutput[41]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U4 ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[40]), .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n13), .A2(AddRoundKeyOutput[43]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n12), .A2(AddRoundKeyOutput[42]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U1 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[24])
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U4 ( .A1(AddRoundKeyOutput[46]), 
        .A2(AddRoundKeyOutput[47]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U3 ( .A1(AddRoundKeyOutput[44]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U2 ( .A1(AddRoundKeyOutput[46]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput[45]), 
        .B(AddRoundKeyOutput[47]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_11_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[25])
         );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(AddRoundKeyOutput[47]), 
        .A2(AddRoundKeyOutput[46]), .ZN(Red_SubCellInst_LFInst_11_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U1 ( .A1(AddRoundKeyOutput[45]), 
        .A2(AddRoundKeyOutput[47]), .ZN(Red_SubCellInst_LFInst_11_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U7 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n17), .A2(
        Red_SubCellInst_LFInst_11_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[26])
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n15), .A2(AddRoundKeyOutput[47]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n14), .A2(AddRoundKeyOutput[46]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U4 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n13), .A2(
        Red_SubCellInst_LFInst_11_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_2_n17) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_2_U2 ( .A(AddRoundKeyOutput[45]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[46]), .Z(Red_SubCellInst_LFInst_11_LFInst_2_n13)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[36])
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U4 ( .A1(AddRoundKeyOutput[50]), 
        .A2(AddRoundKeyOutput[51]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U3 ( .A1(AddRoundKeyOutput[48]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U2 ( .A1(AddRoundKeyOutput[50]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput[49]), 
        .B(AddRoundKeyOutput[51]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_12_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[37])
         );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U2 ( .A1(AddRoundKeyOutput[51]), 
        .A2(AddRoundKeyOutput[50]), .ZN(Red_SubCellInst_LFInst_12_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U1 ( .A1(AddRoundKeyOutput[49]), 
        .A2(AddRoundKeyOutput[51]), .ZN(Red_SubCellInst_LFInst_12_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n16), .A2(
        Red_SubCellInst_LFInst_12_LFInst_2_n15), .ZN(Red_ShiftRowsOutput[38])
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n14), .A2(AddRoundKeyOutput[51]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U4 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n13), .A2(AddRoundKeyOutput[50]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U3 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n13) );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U2 ( .A1(AddRoundKeyOutput[49]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U1 ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[48]), .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[39])
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U4 ( .A1(AddRoundKeyOutput[54]), 
        .A2(AddRoundKeyOutput[55]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U2 ( .A1(AddRoundKeyOutput[54]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput[53]), 
        .B(AddRoundKeyOutput[55]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_13_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[40])
         );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U2 ( .A1(AddRoundKeyOutput[55]), 
        .A2(AddRoundKeyOutput[54]), .ZN(Red_SubCellInst_LFInst_13_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U1 ( .A1(AddRoundKeyOutput[53]), 
        .A2(AddRoundKeyOutput[55]), .ZN(Red_SubCellInst_LFInst_13_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n16), .A2(
        Red_SubCellInst_LFInst_13_LFInst_2_n15), .ZN(Red_ShiftRowsOutput[41])
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n14), .A2(AddRoundKeyOutput[55]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U4 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n13), .A2(AddRoundKeyOutput[54]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n13) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U2 ( .A1(AddRoundKeyOutput[53]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[52]), .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[42])
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U4 ( .A1(AddRoundKeyOutput[58]), 
        .A2(AddRoundKeyOutput[59]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U3 ( .A1(AddRoundKeyOutput[56]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U2 ( .A1(AddRoundKeyOutput[58]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput[57]), 
        .B(AddRoundKeyOutput[59]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_14_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[43])
         );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U2 ( .A1(AddRoundKeyOutput[59]), 
        .A2(AddRoundKeyOutput[58]), .ZN(Red_SubCellInst_LFInst_14_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U1 ( .A1(AddRoundKeyOutput[57]), 
        .A2(AddRoundKeyOutput[59]), .ZN(Red_SubCellInst_LFInst_14_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_14_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[44])
         );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U5 ( .A1(AddRoundKeyOutput[57]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U4 ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[56]), .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n13), .A2(AddRoundKeyOutput[59]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n12), .A2(AddRoundKeyOutput[58]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U1 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[45])
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U4 ( .A1(AddRoundKeyOutput[62]), 
        .A2(AddRoundKeyOutput[63]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U3 ( .A1(AddRoundKeyOutput[60]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U2 ( .A1(AddRoundKeyOutput[62]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput[61]), 
        .B(AddRoundKeyOutput[63]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_15_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[46])
         );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U2 ( .A1(AddRoundKeyOutput[63]), 
        .A2(AddRoundKeyOutput[62]), .ZN(Red_SubCellInst_LFInst_15_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U1 ( .A1(AddRoundKeyOutput[61]), 
        .A2(AddRoundKeyOutput[63]), .ZN(Red_SubCellInst_LFInst_15_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_15_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[47])
         );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U5 ( .A1(AddRoundKeyOutput[61]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U4 ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[60]), .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n13), .A2(AddRoundKeyOutput[63]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n12), .A2(AddRoundKeyOutput[62]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U1 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n12) );
  BUF_X1 Red_MCInst_MC0_U3 ( .A(ShiftRowsOutput[28]), .Z(
        Red_MCInst_MC0_v2_1[1]) );
  BUF_X1 Red_MCInst_MC0_U2 ( .A(MCInst_MC0_v1_3[2]), .Z(Red_MCInst_MC0_v1_2[1]) );
  XOR2_X1 Red_MCInst_MC0_v0_2Inst_0_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(Red_MCInst_MC0_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC0_v0_3Inst_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U2 ( .A(Red_MCInst_MC0_v1_0Inst_0_n3), 
        .B(MCInst_MC0_v1_3[3]), .ZN(Red_MCInst_MC0_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC0_v1_2Inst_0_U1 ( .A(Red_MCInst_MC0_v1_2[1]), .B(
        Red_MCInst_MC0_v1_1[2]), .Z(Red_MCInst_MC0_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC0_v1_3Inst_0_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .Z(Red_MCInst_MC0_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC0_v2_0Inst_0_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(Red_MCInst_MC0_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC0_v2_1Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC0_v2_2Inst_0_U2 ( .A(Red_MCInst_MC0_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC0_v2_2[1]), .ZN(Red_MCInst_MC0_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC0_v2_2Inst_0_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[2]), .ZN(Red_MCInst_MC0_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC0_v2_3Inst_0_U2 ( .A(Red_MCInst_MC0_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC0_v2_2[1]), .ZN(Red_MCInst_MC0_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC0_v2_3Inst_0_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(Red_MCInst_MC0_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC0_v3_0Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U3 ( .A(Red_MCInst_MC0_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC0_v3_2Inst_0_n5), .ZN(Red_MCInst_MC0_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U2 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC0_v3_3Inst_0_U1 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(Red_MCInst_MC0_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC0_v0_0Inst_1_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(Red_MCInst_MC0_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC0_v0_1Inst_1_U2 ( .A(Red_MCInst_MC0_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC0_v0_1[0]), .ZN(Red_MCInst_MC0_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC0_v0_1Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .ZN(Red_MCInst_MC0_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .Z(Red_MCInst_MC0_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_1_U2 ( .A(Red_MCInst_MC0_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_1Inst_1_U3 ( .A(Red_MCInst_MC0_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC0_v1_1Inst_1_n5), .ZN(Red_MCInst_MC0_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC0_v1_1Inst_1_U2 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC0_v1_1Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .Z(Red_MCInst_MC0_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC0_v1_3Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[3]), .Z(Red_MCInst_MC0_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC0_v2_0Inst_1_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC0_v2_3Inst_1_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(Red_MCInst_MC0_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC0_v3_0Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .Z(Red_MCInst_MC0_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC0_v3_1Inst_1_U3 ( .A(Red_MCInst_MC0_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC0_v3_1Inst_1_n5), .ZN(Red_MCInst_MC0_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC0_v3_1Inst_1_U2 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC0_v3_1Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC0_v3_2Inst_1_U1 ( .A(Red_MCInst_MC0_v3_3[2]), .B(
        MCInst_MC0_v3_0[3]), .Z(Red_MCInst_MC0_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC0_v3_3Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC0_v0_0Inst_2_U2 ( .A(Red_MCInst_MC0_v0_0Inst_2_n3), 
        .B(MCInst_MC0_v0_3[3]), .ZN(Red_MCInst_MC0_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .ZN(Red_MCInst_MC0_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC0_v0_1Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_2_U3 ( .A(Red_MCInst_MC0_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC0_v0_3Inst_2_n5), .ZN(Red_MCInst_MC0_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_2_U2 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .ZN(Red_MCInst_MC0_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v0_3Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_2_U2 ( .A(Red_MCInst_MC0_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_2_U1 ( .A(Red_MCInst_MC0_v1_2[1]), .B(
        MCInst_MC0_v1_3[3]), .ZN(Red_MCInst_MC0_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_2Inst_2_U2 ( .A(Red_MCInst_MC0_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC0_v1_2Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_2_U3 ( .A(Red_MCInst_MC0_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC0_v1_3Inst_2_n5), .ZN(Red_MCInst_MC0_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_2_U2 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v1_3Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .Z(Red_MCInst_MC0_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_2_U3 ( .A(Red_MCInst_MC0_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC0_v2_0Inst_2_n5), .ZN(Red_MCInst_MC0_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_2_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(Red_MCInst_MC0_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v2_0Inst_2_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(Red_MCInst_MC0_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC0_v2_1Inst_2_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(Red_MCInst_MC0_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC0_v2_2Inst_2_U1 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(Red_MCInst_MC0_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC0_v2_3Inst_2_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_2_U3 ( .A(Red_MCInst_MC0_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC0_v3_0Inst_2_n5), .ZN(Red_MCInst_MC0_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_2_U2 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v3_0Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_2_U2 ( .A(Red_MCInst_MC0_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .ZN(Red_MCInst_MC0_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[45]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_0[0]), 
        .B(Red_MCInst_MC0_v1_0[0]), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), 
        .B(Red_MCInst_MC0_v3_0[0]), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[46]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_0[1]), 
        .B(Red_MCInst_MC0_v1_0[1]), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_0[1]), 
        .B(Red_MCInst_MC0_v3_0[1]), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[47]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_0[2]), 
        .B(Red_MCInst_MC0_v1_0[2]), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_0[2]), 
        .B(Red_MCInst_MC0_v3_0[2]), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[33]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_1[0]), 
        .B(Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_1[0]), 
        .B(Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[34]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_1[1]), 
        .B(Red_MCInst_MC0_v1_1[1]), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_1[1]), 
        .B(Red_MCInst_MC0_v3_1[1]), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[35]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_1[2]), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_1[2]), 
        .B(Red_MCInst_MC0_v3_1[2]), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[21]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_2[0]), 
        .B(Red_MCInst_MC0_v1_2[0]), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_2[0]), 
        .B(Red_MCInst_MC0_v3_2[0]), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[22]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_2[1]), 
        .B(Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_2[1]), 
        .B(Red_MCInst_MC0_v3_2[1]), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[23]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_2[2]), 
        .B(Red_MCInst_MC0_v1_2[2]), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), 
        .B(Red_MCInst_MC0_v3_2[2]), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[9]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_3[0]), 
        .B(Red_MCInst_MC0_v1_3[0]), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_3[0]), 
        .B(Red_MCInst_MC0_v3_3[0]), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[10]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_3[1]), 
        .B(Red_MCInst_MC0_v1_3[1]), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_3[1]), 
        .B(Red_MCInst_MC0_v3_3[1]), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[11]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_3[2]), 
        .B(Red_MCInst_MC0_v1_3[2]), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_3[2]), 
        .B(Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst_MC1_U3 ( .A(MCInst_MC1_v1_3[2]), .Z(Red_MCInst_MC1_v1_2[1]) );
  BUF_X1 Red_MCInst_MC1_U2 ( .A(ShiftRowsOutput[24]), .Z(
        Red_MCInst_MC1_v2_1[1]) );
  XOR2_X1 Red_MCInst_MC1_v0_2Inst_0_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(Red_MCInst_MC1_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC1_v0_3Inst_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U2 ( .A(Red_MCInst_MC1_v1_0Inst_0_n3), 
        .B(MCInst_MC1_v1_3[3]), .ZN(Red_MCInst_MC1_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC1_v1_2Inst_0_U1 ( .A(Red_MCInst_MC1_v1_2[1]), .B(
        Red_MCInst_MC1_v1_1[2]), .Z(Red_MCInst_MC1_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC1_v1_3Inst_0_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .Z(Red_MCInst_MC1_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC1_v2_0Inst_0_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(Red_MCInst_MC1_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC1_v2_1Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC1_v2_2Inst_0_U2 ( .A(Red_MCInst_MC1_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC1_v2_2[1]), .ZN(Red_MCInst_MC1_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC1_v2_2Inst_0_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[2]), .ZN(Red_MCInst_MC1_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC1_v2_3Inst_0_U2 ( .A(Red_MCInst_MC1_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC1_v2_2[1]), .ZN(Red_MCInst_MC1_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC1_v2_3Inst_0_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(Red_MCInst_MC1_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC1_v3_0Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U3 ( .A(Red_MCInst_MC1_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC1_v3_2Inst_0_n5), .ZN(Red_MCInst_MC1_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U2 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC1_v3_3Inst_0_U1 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(Red_MCInst_MC1_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC1_v0_0Inst_1_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(Red_MCInst_MC1_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC1_v0_1Inst_1_U2 ( .A(Red_MCInst_MC1_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC1_v0_1[0]), .ZN(Red_MCInst_MC1_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC1_v0_1Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .ZN(Red_MCInst_MC1_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .Z(Red_MCInst_MC1_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_1_U2 ( .A(Red_MCInst_MC1_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_1Inst_1_U3 ( .A(Red_MCInst_MC1_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC1_v1_1Inst_1_n5), .ZN(Red_MCInst_MC1_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC1_v1_1Inst_1_U2 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC1_v1_1Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .Z(Red_MCInst_MC1_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC1_v1_3Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[3]), .Z(Red_MCInst_MC1_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC1_v2_0Inst_1_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC1_v2_3Inst_1_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(Red_MCInst_MC1_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC1_v3_0Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .Z(Red_MCInst_MC1_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC1_v3_1Inst_1_U3 ( .A(Red_MCInst_MC1_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC1_v3_1Inst_1_n5), .ZN(Red_MCInst_MC1_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC1_v3_1Inst_1_U2 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC1_v3_1Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC1_v3_2Inst_1_U1 ( .A(Red_MCInst_MC1_v3_3[2]), .B(
        MCInst_MC1_v3_0[3]), .Z(Red_MCInst_MC1_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC1_v3_3Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC1_v0_0Inst_2_U2 ( .A(Red_MCInst_MC1_v0_0Inst_2_n3), 
        .B(MCInst_MC1_v0_3[3]), .ZN(Red_MCInst_MC1_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .ZN(Red_MCInst_MC1_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC1_v0_1Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_2_U3 ( .A(Red_MCInst_MC1_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC1_v0_3Inst_2_n5), .ZN(Red_MCInst_MC1_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_2_U2 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .ZN(Red_MCInst_MC1_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v0_3Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_2_U2 ( .A(Red_MCInst_MC1_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_2_U1 ( .A(Red_MCInst_MC1_v1_2[1]), .B(
        MCInst_MC1_v1_3[3]), .ZN(Red_MCInst_MC1_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_2Inst_2_U2 ( .A(Red_MCInst_MC1_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC1_v1_2Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_2_U3 ( .A(Red_MCInst_MC1_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC1_v1_3Inst_2_n5), .ZN(Red_MCInst_MC1_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_2_U2 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v1_3Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .Z(Red_MCInst_MC1_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_2_U3 ( .A(Red_MCInst_MC1_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC1_v2_0Inst_2_n5), .ZN(Red_MCInst_MC1_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_2_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(Red_MCInst_MC1_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v2_0Inst_2_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(Red_MCInst_MC1_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC1_v2_1Inst_2_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(Red_MCInst_MC1_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC1_v2_2Inst_2_U1 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(Red_MCInst_MC1_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC1_v2_3Inst_2_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_2_U3 ( .A(Red_MCInst_MC1_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC1_v3_0Inst_2_n5), .ZN(Red_MCInst_MC1_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_2_U2 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v3_0Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_2_U2 ( .A(Red_MCInst_MC1_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .ZN(Red_MCInst_MC1_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[42]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_0[0]), 
        .B(Red_MCInst_MC1_v1_0[0]), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), 
        .B(Red_MCInst_MC1_v3_0[0]), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[43]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_0[1]), 
        .B(Red_MCInst_MC1_v1_0[1]), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_0[1]), 
        .B(Red_MCInst_MC1_v3_0[1]), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[44]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_0[2]), 
        .B(Red_MCInst_MC1_v1_0[2]), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_0[2]), 
        .B(Red_MCInst_MC1_v3_0[2]), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[30]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_1[0]), 
        .B(Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_1[0]), 
        .B(Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[31]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_1[1]), 
        .B(Red_MCInst_MC1_v1_1[1]), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_1[1]), 
        .B(Red_MCInst_MC1_v3_1[1]), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[32]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_1[2]), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_1[2]), 
        .B(Red_MCInst_MC1_v3_1[2]), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[18]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_2[0]), 
        .B(Red_MCInst_MC1_v1_2[0]), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_2[0]), 
        .B(Red_MCInst_MC1_v3_2[0]), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[19]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_2[1]), 
        .B(Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_2[1]), 
        .B(Red_MCInst_MC1_v3_2[1]), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[20]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_2[2]), 
        .B(Red_MCInst_MC1_v1_2[2]), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), 
        .B(Red_MCInst_MC1_v3_2[2]), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[6]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_3[0]), 
        .B(Red_MCInst_MC1_v1_3[0]), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_3[0]), 
        .B(Red_MCInst_MC1_v3_3[0]), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[7]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_3[1]), 
        .B(Red_MCInst_MC1_v1_3[1]), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_3[1]), 
        .B(Red_MCInst_MC1_v3_3[1]), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[8]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_3[2]), 
        .B(Red_MCInst_MC1_v1_3[2]), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_3[2]), 
        .B(Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst_MC2_U3 ( .A(MCInst_MC2_v1_3[2]), .Z(Red_MCInst_MC2_v1_2[1]) );
  BUF_X1 Red_MCInst_MC2_U2 ( .A(ShiftRowsOutput[20]), .Z(
        Red_MCInst_MC2_v2_1[1]) );
  XOR2_X1 Red_MCInst_MC2_v0_2Inst_0_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(Red_MCInst_MC2_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC2_v0_3Inst_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U2 ( .A(Red_MCInst_MC2_v1_0Inst_0_n3), 
        .B(MCInst_MC2_v1_3[3]), .ZN(Red_MCInst_MC2_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC2_v1_2Inst_0_U1 ( .A(Red_MCInst_MC2_v1_2[1]), .B(
        Red_MCInst_MC2_v1_1[2]), .Z(Red_MCInst_MC2_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC2_v1_3Inst_0_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .Z(Red_MCInst_MC2_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC2_v2_0Inst_0_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(Red_MCInst_MC2_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC2_v2_1Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC2_v2_2Inst_0_U2 ( .A(Red_MCInst_MC2_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC2_v2_2[1]), .ZN(Red_MCInst_MC2_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC2_v2_2Inst_0_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[2]), .ZN(Red_MCInst_MC2_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC2_v2_3Inst_0_U2 ( .A(Red_MCInst_MC2_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC2_v2_2[1]), .ZN(Red_MCInst_MC2_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC2_v2_3Inst_0_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(Red_MCInst_MC2_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC2_v3_0Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U3 ( .A(Red_MCInst_MC2_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC2_v3_2Inst_0_n5), .ZN(Red_MCInst_MC2_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U2 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC2_v3_3Inst_0_U1 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(Red_MCInst_MC2_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC2_v0_0Inst_1_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(Red_MCInst_MC2_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC2_v0_1Inst_1_U2 ( .A(Red_MCInst_MC2_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC2_v0_1[0]), .ZN(Red_MCInst_MC2_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC2_v0_1Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .ZN(Red_MCInst_MC2_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .Z(Red_MCInst_MC2_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_1_U2 ( .A(Red_MCInst_MC2_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_1Inst_1_U3 ( .A(Red_MCInst_MC2_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC2_v1_1Inst_1_n5), .ZN(Red_MCInst_MC2_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC2_v1_1Inst_1_U2 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC2_v1_1Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .Z(Red_MCInst_MC2_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC2_v1_3Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[3]), .Z(Red_MCInst_MC2_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC2_v2_0Inst_1_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC2_v2_3Inst_1_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(Red_MCInst_MC2_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC2_v3_0Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .Z(Red_MCInst_MC2_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC2_v3_1Inst_1_U3 ( .A(Red_MCInst_MC2_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC2_v3_1Inst_1_n5), .ZN(Red_MCInst_MC2_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC2_v3_1Inst_1_U2 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC2_v3_1Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC2_v3_2Inst_1_U1 ( .A(Red_MCInst_MC2_v3_3[2]), .B(
        MCInst_MC2_v3_0[3]), .Z(Red_MCInst_MC2_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC2_v3_3Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC2_v0_0Inst_2_U2 ( .A(Red_MCInst_MC2_v0_0Inst_2_n3), 
        .B(MCInst_MC2_v0_3[3]), .ZN(Red_MCInst_MC2_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .ZN(Red_MCInst_MC2_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC2_v0_1Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_2_U3 ( .A(Red_MCInst_MC2_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC2_v0_3Inst_2_n5), .ZN(Red_MCInst_MC2_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_2_U2 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .ZN(Red_MCInst_MC2_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v0_3Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_2_U2 ( .A(Red_MCInst_MC2_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_2_U1 ( .A(Red_MCInst_MC2_v1_2[1]), .B(
        MCInst_MC2_v1_3[3]), .ZN(Red_MCInst_MC2_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_2Inst_2_U2 ( .A(Red_MCInst_MC2_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC2_v1_2Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_2_U3 ( .A(Red_MCInst_MC2_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC2_v1_3Inst_2_n5), .ZN(Red_MCInst_MC2_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_2_U2 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v1_3Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .Z(Red_MCInst_MC2_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_2_U3 ( .A(Red_MCInst_MC2_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC2_v2_0Inst_2_n5), .ZN(Red_MCInst_MC2_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_2_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(Red_MCInst_MC2_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v2_0Inst_2_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(Red_MCInst_MC2_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC2_v2_1Inst_2_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(Red_MCInst_MC2_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC2_v2_2Inst_2_U1 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(Red_MCInst_MC2_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC2_v2_3Inst_2_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_2_U3 ( .A(Red_MCInst_MC2_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC2_v3_0Inst_2_n5), .ZN(Red_MCInst_MC2_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_2_U2 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v3_0Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_2_U2 ( .A(Red_MCInst_MC2_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .ZN(Red_MCInst_MC2_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[39]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_0[0]), 
        .B(Red_MCInst_MC2_v1_0[0]), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), 
        .B(Red_MCInst_MC2_v3_0[0]), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[40]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_0[1]), 
        .B(Red_MCInst_MC2_v1_0[1]), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_0[1]), 
        .B(Red_MCInst_MC2_v3_0[1]), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[41]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_0[2]), 
        .B(Red_MCInst_MC2_v1_0[2]), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_0[2]), 
        .B(Red_MCInst_MC2_v3_0[2]), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[27]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_1[0]), 
        .B(Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_1[0]), 
        .B(Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[28]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_1[1]), 
        .B(Red_MCInst_MC2_v1_1[1]), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_1[1]), 
        .B(Red_MCInst_MC2_v3_1[1]), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[29]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_1[2]), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_1[2]), 
        .B(Red_MCInst_MC2_v3_1[2]), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[15]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_2[0]), 
        .B(Red_MCInst_MC2_v1_2[0]), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_2[0]), 
        .B(Red_MCInst_MC2_v3_2[0]), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[16]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_2[1]), 
        .B(Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_2[1]), 
        .B(Red_MCInst_MC2_v3_2[1]), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[17]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_2[2]), 
        .B(Red_MCInst_MC2_v1_2[2]), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), 
        .B(Red_MCInst_MC2_v3_2[2]), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[3]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_3[0]), 
        .B(Red_MCInst_MC2_v1_3[0]), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_3[0]), 
        .B(Red_MCInst_MC2_v3_3[0]), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[4]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_3[1]), 
        .B(Red_MCInst_MC2_v1_3[1]), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_3[1]), 
        .B(Red_MCInst_MC2_v3_3[1]), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[5]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_3[2]), 
        .B(Red_MCInst_MC2_v1_3[2]), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_3[2]), 
        .B(Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst_MC3_U3 ( .A(ShiftRowsOutput[16]), .Z(
        Red_MCInst_MC3_v2_1[1]) );
  BUF_X1 Red_MCInst_MC3_U2 ( .A(MCInst_MC3_v1_3[2]), .Z(Red_MCInst_MC3_v1_2[1]) );
  XOR2_X1 Red_MCInst_MC3_v0_2Inst_0_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(Red_MCInst_MC3_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC3_v0_3Inst_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U2 ( .A(Red_MCInst_MC3_v1_0Inst_0_n3), 
        .B(MCInst_MC3_v1_3[3]), .ZN(Red_MCInst_MC3_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC3_v1_2Inst_0_U1 ( .A(Red_MCInst_MC3_v1_2[1]), .B(
        Red_MCInst_MC3_v1_1[2]), .Z(Red_MCInst_MC3_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC3_v1_3Inst_0_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .Z(Red_MCInst_MC3_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC3_v2_0Inst_0_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(Red_MCInst_MC3_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC3_v2_1Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC3_v2_2Inst_0_U2 ( .A(Red_MCInst_MC3_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC3_v2_2[1]), .ZN(Red_MCInst_MC3_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC3_v2_2Inst_0_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[2]), .ZN(Red_MCInst_MC3_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC3_v2_3Inst_0_U2 ( .A(Red_MCInst_MC3_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC3_v2_2[1]), .ZN(Red_MCInst_MC3_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC3_v2_3Inst_0_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(Red_MCInst_MC3_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC3_v3_0Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U3 ( .A(Red_MCInst_MC3_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC3_v3_2Inst_0_n5), .ZN(Red_MCInst_MC3_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U2 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC3_v3_3Inst_0_U1 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(Red_MCInst_MC3_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC3_v0_0Inst_1_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(Red_MCInst_MC3_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC3_v0_1Inst_1_U2 ( .A(Red_MCInst_MC3_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC3_v0_1[0]), .ZN(Red_MCInst_MC3_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC3_v0_1Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .ZN(Red_MCInst_MC3_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .Z(Red_MCInst_MC3_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_1_U2 ( .A(Red_MCInst_MC3_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_1Inst_1_U3 ( .A(Red_MCInst_MC3_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC3_v1_1Inst_1_n5), .ZN(Red_MCInst_MC3_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC3_v1_1Inst_1_U2 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC3_v1_1Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .Z(Red_MCInst_MC3_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC3_v1_3Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[3]), .Z(Red_MCInst_MC3_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC3_v2_0Inst_1_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC3_v2_3Inst_1_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(Red_MCInst_MC3_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC3_v3_0Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .Z(Red_MCInst_MC3_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC3_v3_1Inst_1_U3 ( .A(Red_MCInst_MC3_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC3_v3_1Inst_1_n5), .ZN(Red_MCInst_MC3_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC3_v3_1Inst_1_U2 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC3_v3_1Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC3_v3_2Inst_1_U1 ( .A(Red_MCInst_MC3_v3_3[2]), .B(
        MCInst_MC3_v3_0[3]), .Z(Red_MCInst_MC3_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC3_v3_3Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC3_v0_0Inst_2_U2 ( .A(Red_MCInst_MC3_v0_0Inst_2_n3), 
        .B(MCInst_MC3_v0_3[3]), .ZN(Red_MCInst_MC3_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .ZN(Red_MCInst_MC3_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC3_v0_1Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_2_U3 ( .A(Red_MCInst_MC3_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC3_v0_3Inst_2_n5), .ZN(Red_MCInst_MC3_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_2_U2 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .ZN(Red_MCInst_MC3_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v0_3Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_2_U2 ( .A(Red_MCInst_MC3_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_2_U1 ( .A(Red_MCInst_MC3_v1_2[1]), .B(
        MCInst_MC3_v1_3[3]), .ZN(Red_MCInst_MC3_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_2Inst_2_U2 ( .A(Red_MCInst_MC3_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC3_v1_2Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_2_U3 ( .A(Red_MCInst_MC3_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC3_v1_3Inst_2_n5), .ZN(Red_MCInst_MC3_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_2_U2 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v1_3Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .Z(Red_MCInst_MC3_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_2_U3 ( .A(Red_MCInst_MC3_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC3_v2_0Inst_2_n5), .ZN(Red_MCInst_MC3_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_2_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(Red_MCInst_MC3_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v2_0Inst_2_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(Red_MCInst_MC3_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC3_v2_1Inst_2_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(Red_MCInst_MC3_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC3_v2_2Inst_2_U1 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(Red_MCInst_MC3_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC3_v2_3Inst_2_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_2_U3 ( .A(Red_MCInst_MC3_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC3_v3_0Inst_2_n5), .ZN(Red_MCInst_MC3_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_2_U2 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v3_0Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_2_U2 ( .A(Red_MCInst_MC3_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .ZN(Red_MCInst_MC3_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[36]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_0[0]), 
        .B(Red_MCInst_MC3_v1_0[0]), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), 
        .B(Red_MCInst_MC3_v3_0[0]), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[37]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_0[1]), 
        .B(Red_MCInst_MC3_v1_0[1]), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_0[1]), 
        .B(Red_MCInst_MC3_v3_0[1]), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[38]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_0[2]), 
        .B(Red_MCInst_MC3_v1_0[2]), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_0[2]), 
        .B(Red_MCInst_MC3_v3_0[2]), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[24]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_1[0]), 
        .B(Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_1[0]), 
        .B(Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[25]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_1[1]), 
        .B(Red_MCInst_MC3_v1_1[1]), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_1[1]), 
        .B(Red_MCInst_MC3_v3_1[1]), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[26]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_1[2]), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_1[2]), 
        .B(Red_MCInst_MC3_v3_1[2]), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[12]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_2[0]), 
        .B(Red_MCInst_MC3_v1_2[0]), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_2[0]), 
        .B(Red_MCInst_MC3_v3_2[0]), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[13]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_2[1]), 
        .B(Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_2[1]), 
        .B(Red_MCInst_MC3_v3_2[1]), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[14]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_2[2]), 
        .B(Red_MCInst_MC3_v1_2[2]), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), 
        .B(Red_MCInst_MC3_v3_2[2]), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[0]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_3[0]), 
        .B(Red_MCInst_MC3_v1_3[0]), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_3[0]), 
        .B(Red_MCInst_MC3_v3_3[0]), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[1]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_3[1]), 
        .B(Red_MCInst_MC3_v1_3[1]), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_3[1]), 
        .B(Red_MCInst_MC3_v3_3[1]), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[2]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_3[2]), 
        .B(Red_MCInst_MC3_v1_3[2]), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_3[2]), 
        .B(Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_0_LFInst_0_n3), .B(Key[2]), .ZN(Red_RoundKey[0]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_0_LFInst_1_n3), .B(Key[3]), .ZN(Red_RoundKey[1]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_1_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_0_LFInst_2_n3), .B(Key[3]), .ZN(Red_RoundKey[2]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_2_U1 ( .A(Key[1]), .B(Key[2]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_1_LFInst_0_n3), .B(Key[6]), .ZN(Red_RoundKey[3]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_1_LFInst_1_n3), .B(Key[7]), .ZN(Red_RoundKey[4]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_1_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_1_LFInst_2_n3), .B(Key[7]), .ZN(Red_RoundKey[5]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_2_U1 ( .A(Key[5]), .B(Key[6]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_2_LFInst_0_n3), .B(Key[10]), .ZN(Red_RoundKey[6])
         );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_2_LFInst_1_n3), .B(Key[11]), .ZN(Red_RoundKey[7])
         );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_1_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_2_LFInst_2_n3), .B(Key[11]), .ZN(Red_RoundKey[8])
         );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_2_U1 ( .A(Key[9]), .B(Key[10]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_3_LFInst_0_n3), .B(Key[14]), .ZN(Red_RoundKey[9])
         );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_3_LFInst_1_n3), .B(Key[15]), .ZN(Red_RoundKey[10])
         );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_1_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_3_LFInst_2_n3), .B(Key[15]), .ZN(Red_RoundKey[11])
         );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_2_U1 ( .A(Key[13]), .B(Key[14]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_4_LFInst_0_n3), .B(Key[18]), .ZN(Red_RoundKey[12])
         );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_4_LFInst_1_n3), .B(Key[19]), .ZN(Red_RoundKey[13])
         );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_1_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_4_LFInst_2_n3), .B(Key[19]), .ZN(Red_RoundKey[14])
         );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_2_U1 ( .A(Key[17]), .B(Key[18]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_5_LFInst_0_n3), .B(Key[22]), .ZN(Red_RoundKey[15])
         );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_5_LFInst_1_n3), .B(Key[23]), .ZN(Red_RoundKey[16])
         );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_1_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_5_LFInst_2_n3), .B(Key[23]), .ZN(Red_RoundKey[17])
         );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_2_U1 ( .A(Key[21]), .B(Key[22]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_6_LFInst_0_n3), .B(Key[26]), .ZN(Red_RoundKey[18])
         );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_6_LFInst_1_n3), .B(Key[27]), .ZN(Red_RoundKey[19])
         );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_1_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_6_LFInst_2_n3), .B(Key[27]), .ZN(Red_RoundKey[20])
         );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_2_U1 ( .A(Key[25]), .B(Key[26]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_7_LFInst_0_n3), .B(Key[30]), .ZN(Red_RoundKey[21])
         );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_7_LFInst_1_n3), .B(Key[31]), .ZN(Red_RoundKey[22])
         );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_1_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_7_LFInst_2_n3), .B(Key[31]), .ZN(Red_RoundKey[23])
         );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_2_U1 ( .A(Key[29]), .B(Key[30]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_8_LFInst_0_n3), .B(Key[34]), .ZN(Red_RoundKey[24])
         );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_8_LFInst_1_n3), .B(Key[35]), .ZN(Red_RoundKey[25])
         );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_1_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_8_LFInst_2_n3), .B(Key[35]), .ZN(Red_RoundKey[26])
         );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_2_U1 ( .A(Key[33]), .B(Key[34]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_9_LFInst_0_n3), .B(Key[38]), .ZN(Red_RoundKey[27])
         );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_9_LFInst_1_n3), .B(Key[39]), .ZN(Red_RoundKey[28])
         );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_1_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_9_LFInst_2_n3), .B(Key[39]), .ZN(Red_RoundKey[29])
         );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_2_U1 ( .A(Key[37]), .B(Key[38]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_10_LFInst_0_n3), .B(Key[42]), .ZN(Red_RoundKey[30])
         );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_10_LFInst_1_n3), .B(Key[43]), .ZN(Red_RoundKey[31])
         );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_1_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_10_LFInst_2_n3), .B(Key[43]), .ZN(Red_RoundKey[32])
         );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_2_U1 ( .A(Key[41]), .B(Key[42]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_11_LFInst_0_n3), .B(Key[46]), .ZN(Red_RoundKey[33])
         );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_11_LFInst_1_n3), .B(Key[47]), .ZN(Red_RoundKey[34])
         );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_1_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_11_LFInst_2_n3), .B(Key[47]), .ZN(Red_RoundKey[35])
         );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_2_U1 ( .A(Key[45]), .B(Key[46]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_12_LFInst_0_n3), .B(Key[50]), .ZN(Red_RoundKey[36])
         );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_12_LFInst_1_n3), .B(Key[51]), .ZN(Red_RoundKey[37])
         );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_1_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_12_LFInst_2_n3), .B(Key[51]), .ZN(Red_RoundKey[38])
         );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_2_U1 ( .A(Key[49]), .B(Key[50]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_13_LFInst_0_n3), .B(Key[54]), .ZN(Red_RoundKey[39])
         );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_13_LFInst_1_n3), .B(Key[55]), .ZN(Red_RoundKey[40])
         );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_1_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_13_LFInst_2_n3), .B(Key[55]), .ZN(Red_RoundKey[41])
         );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_2_U1 ( .A(Key[53]), .B(Key[54]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_14_LFInst_0_n3), .B(Key[58]), .ZN(Red_RoundKey[42])
         );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_14_LFInst_1_n3), .B(Key[59]), .ZN(Red_RoundKey[43])
         );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_1_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_14_LFInst_2_n3), .B(Key[59]), .ZN(Red_RoundKey[44])
         );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_2_U1 ( .A(Key[57]), .B(Key[58]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_15_LFInst_0_n3), .B(Key[62]), .ZN(Red_RoundKey[45])
         );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_15_LFInst_1_n3), .B(Key[63]), .ZN(Red_RoundKey[46])
         );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_1_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_15_LFInst_2_n3), .B(Key[63]), .ZN(Red_RoundKey[47])
         );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_2_U1 ( .A(Key[61]), .B(Key[62]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_0_n3), .B(AddRoundKeyOutput[2]), .ZN(
        Red_SignaltoCheck[0]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_1_n3), .B(AddRoundKeyOutput[3]), .ZN(
        Red_SignaltoCheck[1]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_1_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_2_n3), .B(AddRoundKeyOutput[3]), .ZN(
        Red_SignaltoCheck[2]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[1]), 
        .B(AddRoundKeyOutput[2]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_0_n3), .B(AddRoundKeyOutput[6]), .ZN(
        Red_SignaltoCheck[3]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_1_n3), .B(AddRoundKeyOutput[7]), .ZN(
        Red_SignaltoCheck[4]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_1_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_2_n3), .B(AddRoundKeyOutput[7]), .ZN(
        Red_SignaltoCheck[5]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[5]), 
        .B(AddRoundKeyOutput[6]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_0_n3), .B(AddRoundKeyOutput[10]), .ZN(
        Red_SignaltoCheck[6]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_1_n3), .B(AddRoundKeyOutput[11]), .ZN(
        Red_SignaltoCheck[7]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_1_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_2_n3), .B(AddRoundKeyOutput[11]), .ZN(
        Red_SignaltoCheck[8]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_2_U1 ( .A(AddRoundKeyOutput[9]), 
        .B(AddRoundKeyOutput[10]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_0_n3), .B(AddRoundKeyOutput[14]), .ZN(
        Red_SignaltoCheck[9]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_1_n3), .B(AddRoundKeyOutput[15]), .ZN(
        Red_SignaltoCheck[10]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_1_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_2_n3), .B(AddRoundKeyOutput[15]), .ZN(
        Red_SignaltoCheck[11]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_2_U1 ( .A(AddRoundKeyOutput[13]), 
        .B(AddRoundKeyOutput[14]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_0_n3), .B(AddRoundKeyOutput[18]), .ZN(
        Red_SignaltoCheck[12]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_1_n3), .B(AddRoundKeyOutput[19]), .ZN(
        Red_SignaltoCheck[13]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_1_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_2_n3), .B(AddRoundKeyOutput[19]), .ZN(
        Red_SignaltoCheck[14]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_2_U1 ( .A(AddRoundKeyOutput[17]), 
        .B(AddRoundKeyOutput[18]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_0_n3), .B(AddRoundKeyOutput[22]), .ZN(
        Red_SignaltoCheck[15]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_1_n3), .B(AddRoundKeyOutput[23]), .ZN(
        Red_SignaltoCheck[16]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_1_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_2_n3), .B(AddRoundKeyOutput[23]), .ZN(
        Red_SignaltoCheck[17]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_2_U1 ( .A(AddRoundKeyOutput[21]), 
        .B(AddRoundKeyOutput[22]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_0_n3), .B(AddRoundKeyOutput[26]), .ZN(
        Red_SignaltoCheck[18]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_1_n3), .B(AddRoundKeyOutput[27]), .ZN(
        Red_SignaltoCheck[19]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_1_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_2_n3), .B(AddRoundKeyOutput[27]), .ZN(
        Red_SignaltoCheck[20]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_2_U1 ( .A(AddRoundKeyOutput[25]), 
        .B(AddRoundKeyOutput[26]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_0_n3), .B(AddRoundKeyOutput[30]), .ZN(
        Red_SignaltoCheck[21]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_1_n3), .B(AddRoundKeyOutput[31]), .ZN(
        Red_SignaltoCheck[22]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_1_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_2_n3), .B(AddRoundKeyOutput[31]), .ZN(
        Red_SignaltoCheck[23]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_2_U1 ( .A(AddRoundKeyOutput[29]), 
        .B(AddRoundKeyOutput[30]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_0_n3), .B(AddRoundKeyOutput[34]), .ZN(
        Red_SignaltoCheck[24]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_1_n3), .B(AddRoundKeyOutput[35]), .ZN(
        Red_SignaltoCheck[25]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_1_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_2_n3), .B(AddRoundKeyOutput[35]), .ZN(
        Red_SignaltoCheck[26]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_2_U1 ( .A(AddRoundKeyOutput[33]), 
        .B(AddRoundKeyOutput[34]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_0_n3), .B(AddRoundKeyOutput[38]), .ZN(
        Red_SignaltoCheck[27]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_1_n3), .B(AddRoundKeyOutput[39]), .ZN(
        Red_SignaltoCheck[28]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_1_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_2_n3), .B(AddRoundKeyOutput[39]), .ZN(
        Red_SignaltoCheck[29]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_2_U1 ( .A(AddRoundKeyOutput[37]), 
        .B(AddRoundKeyOutput[38]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_0_n3), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_1_n3), .B(AddRoundKeyOutput[43]), 
        .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_1_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_2_n3), .B(AddRoundKeyOutput[43]), 
        .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_2_U1 ( .A(AddRoundKeyOutput[41]), 
        .B(AddRoundKeyOutput[42]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_0_n3), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_1_n3), .B(AddRoundKeyOutput[47]), 
        .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_1_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_2_n3), .B(AddRoundKeyOutput[47]), 
        .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[45]), 
        .B(AddRoundKeyOutput[46]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_0_n3), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_1_n3), .B(AddRoundKeyOutput[51]), 
        .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_1_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_2_n3), .B(AddRoundKeyOutput[51]), 
        .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_2_U1 ( .A(AddRoundKeyOutput[49]), 
        .B(AddRoundKeyOutput[50]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_0_n3), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_1_n3), .B(AddRoundKeyOutput[55]), 
        .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_1_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_2_n3), .B(AddRoundKeyOutput[55]), 
        .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[53]), 
        .B(AddRoundKeyOutput[54]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_0_n3), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_1_n3), .B(AddRoundKeyOutput[59]), 
        .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_1_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_2_n3), .B(AddRoundKeyOutput[59]), 
        .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_2_U1 ( .A(AddRoundKeyOutput[57]), 
        .B(AddRoundKeyOutput[58]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_0_n3), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_1_n3), .B(AddRoundKeyOutput[63]), 
        .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_1_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_2_n3), .B(AddRoundKeyOutput[63]), 
        .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_2_U1 ( .A(AddRoundKeyOutput[61]), 
        .B(AddRoundKeyOutput[62]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_0_n3), .B(Ciphertext[2]), .ZN(
        Red_SignaltoCheck[48]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U1 ( .A(Ciphertext[0]), .B(
        Ciphertext[1]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_1_n3), .B(Ciphertext[3]), .ZN(
        Red_SignaltoCheck[49]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_1_U1 ( .A(Ciphertext[0]), .B(
        Ciphertext[1]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_2_n3), .B(Ciphertext[3]), .ZN(
        Red_SignaltoCheck[50]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_2_U1 ( .A(Ciphertext[1]), .B(
        Ciphertext[2]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_0_n3), .B(Ciphertext[6]), .ZN(
        Red_SignaltoCheck[51]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U1 ( .A(Ciphertext[4]), .B(
        Ciphertext[5]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_1_n3), .B(Ciphertext[7]), .ZN(
        Red_SignaltoCheck[52]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_1_U1 ( .A(Ciphertext[4]), .B(
        Ciphertext[5]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_2_n3), .B(Ciphertext[7]), .ZN(
        Red_SignaltoCheck[53]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_2_U1 ( .A(Ciphertext[5]), .B(
        Ciphertext[6]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_0_n3), .B(Ciphertext[10]), .ZN(
        Red_SignaltoCheck[54]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U1 ( .A(Ciphertext[8]), .B(
        Ciphertext[9]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_1_n3), .B(Ciphertext[11]), .ZN(
        Red_SignaltoCheck[55]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_1_U1 ( .A(Ciphertext[8]), .B(
        Ciphertext[9]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_2_n3), .B(Ciphertext[11]), .ZN(
        Red_SignaltoCheck[56]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_2_U1 ( .A(Ciphertext[9]), .B(
        Ciphertext[10]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_0_n3), .B(Ciphertext[14]), .ZN(
        Red_SignaltoCheck[57]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U1 ( .A(Ciphertext[12]), .B(
        Ciphertext[13]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_1_n3), .B(Ciphertext[15]), .ZN(
        Red_SignaltoCheck[58]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_1_U1 ( .A(Ciphertext[12]), .B(
        Ciphertext[13]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_2_n3), .B(Ciphertext[15]), .ZN(
        Red_SignaltoCheck[59]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_2_U1 ( .A(Ciphertext[13]), .B(
        Ciphertext[14]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_0_n3), .B(Ciphertext[18]), .ZN(
        Red_SignaltoCheck[60]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U1 ( .A(Ciphertext[16]), .B(
        Ciphertext[17]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_1_n3), .B(Ciphertext[19]), .ZN(
        Red_SignaltoCheck[61]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_1_U1 ( .A(Ciphertext[16]), .B(
        Ciphertext[17]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_2_n3), .B(Ciphertext[19]), .ZN(
        Red_SignaltoCheck[62]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_2_U1 ( .A(Ciphertext[17]), .B(
        Ciphertext[18]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_0_n3), .B(Ciphertext[22]), .ZN(
        Red_SignaltoCheck[63]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U1 ( .A(Ciphertext[20]), .B(
        Ciphertext[21]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_1_n3), .B(Ciphertext[23]), .ZN(
        Red_SignaltoCheck[64]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_1_U1 ( .A(Ciphertext[20]), .B(
        Ciphertext[21]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_2_n3), .B(Ciphertext[23]), .ZN(
        Red_SignaltoCheck[65]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_2_U1 ( .A(Ciphertext[21]), .B(
        Ciphertext[22]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_0_n3), .B(Ciphertext[26]), .ZN(
        Red_SignaltoCheck[66]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U1 ( .A(Ciphertext[24]), .B(
        Ciphertext[25]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_1_n3), .B(Ciphertext[27]), .ZN(
        Red_SignaltoCheck[67]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_1_U1 ( .A(Ciphertext[24]), .B(
        Ciphertext[25]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_2_n3), .B(Ciphertext[27]), .ZN(
        Red_SignaltoCheck[68]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_2_U1 ( .A(Ciphertext[25]), .B(
        Ciphertext[26]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_0_n3), .B(Ciphertext[30]), .ZN(
        Red_SignaltoCheck[69]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U1 ( .A(Ciphertext[28]), .B(
        Ciphertext[29]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_1_n3), .B(Ciphertext[31]), .ZN(
        Red_SignaltoCheck[70]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_1_U1 ( .A(Ciphertext[28]), .B(
        Ciphertext[29]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_2_n3), .B(Ciphertext[31]), .ZN(
        Red_SignaltoCheck[71]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_2_U1 ( .A(Ciphertext[29]), .B(
        Ciphertext[30]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_0_n3), .B(Ciphertext[34]), .ZN(
        Red_SignaltoCheck[72]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U1 ( .A(Ciphertext[32]), .B(
        Ciphertext[33]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_1_n3), .B(Ciphertext[35]), .ZN(
        Red_SignaltoCheck[73]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_1_U1 ( .A(Ciphertext[32]), .B(
        Ciphertext[33]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_2_n3), .B(Ciphertext[35]), .ZN(
        Red_SignaltoCheck[74]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_2_U1 ( .A(Ciphertext[33]), .B(
        Ciphertext[34]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_0_n3), .B(Ciphertext[38]), .ZN(
        Red_SignaltoCheck[75]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U1 ( .A(Ciphertext[36]), .B(
        Ciphertext[37]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_1_n3), .B(Ciphertext[39]), .ZN(
        Red_SignaltoCheck[76]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_1_U1 ( .A(Ciphertext[36]), .B(
        Ciphertext[37]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_2_n3), .B(Ciphertext[39]), .ZN(
        Red_SignaltoCheck[77]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_2_U1 ( .A(Ciphertext[37]), .B(
        Ciphertext[38]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_0_n3), .B(Ciphertext[42]), .ZN(
        Red_SignaltoCheck[78]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U1 ( .A(Ciphertext[40]), .B(
        Ciphertext[41]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_1_n3), .B(Ciphertext[43]), .ZN(
        Red_SignaltoCheck[79]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_1_U1 ( .A(Ciphertext[40]), .B(
        Ciphertext[41]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_2_n3), .B(Ciphertext[43]), .ZN(
        Red_SignaltoCheck[80]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_2_U1 ( .A(Ciphertext[41]), .B(
        Ciphertext[42]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_0_n3), .B(Ciphertext[46]), .ZN(
        Red_SignaltoCheck[81]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U1 ( .A(Ciphertext[44]), .B(
        Ciphertext[45]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_1_n3), .B(Ciphertext[47]), .ZN(
        Red_SignaltoCheck[82]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_1_U1 ( .A(Ciphertext[44]), .B(
        Ciphertext[45]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_2_n3), .B(Ciphertext[47]), .ZN(
        Red_SignaltoCheck[83]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_2_U1 ( .A(Ciphertext[45]), .B(
        Ciphertext[46]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_0_n3), .B(Ciphertext[50]), .ZN(
        Red_SignaltoCheck[84]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U1 ( .A(Ciphertext[48]), .B(
        Ciphertext[49]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_1_n3), .B(Ciphertext[51]), .ZN(
        Red_SignaltoCheck[85]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_1_U1 ( .A(Ciphertext[48]), .B(
        Ciphertext[49]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_2_n3), .B(Ciphertext[51]), .ZN(
        Red_SignaltoCheck[86]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_2_U1 ( .A(Ciphertext[49]), .B(
        Ciphertext[50]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_0_n3), .B(Ciphertext[54]), .ZN(
        Red_SignaltoCheck[87]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U1 ( .A(Ciphertext[52]), .B(
        Ciphertext[53]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_1_n3), .B(Ciphertext[55]), .ZN(
        Red_SignaltoCheck[88]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_1_U1 ( .A(Ciphertext[52]), .B(
        Ciphertext[53]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_2_n3), .B(Ciphertext[55]), .ZN(
        Red_SignaltoCheck[89]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_2_U1 ( .A(Ciphertext[53]), .B(
        Ciphertext[54]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_0_n3), .B(Ciphertext[58]), .ZN(
        Red_SignaltoCheck[90]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U1 ( .A(Ciphertext[56]), .B(
        Ciphertext[57]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_1_n3), .B(Ciphertext[59]), .ZN(
        Red_SignaltoCheck[91]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_1_U1 ( .A(Ciphertext[56]), .B(
        Ciphertext[57]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_2_n3), .B(Ciphertext[59]), .ZN(
        Red_SignaltoCheck[92]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_2_U1 ( .A(Ciphertext[57]), .B(
        Ciphertext[58]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_0_n3), .B(Ciphertext[62]), .ZN(
        Red_SignaltoCheck[93]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U1 ( .A(Ciphertext[60]), .B(
        Ciphertext[61]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_1_n3), .B(Ciphertext[63]), .ZN(
        Red_SignaltoCheck[94]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_1_U1 ( .A(Ciphertext[60]), .B(
        Ciphertext[61]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_2_n3), .B(Ciphertext[63]), .ZN(
        Red_SignaltoCheck[95]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_2_U1 ( .A(Ciphertext[61]), .B(
        Ciphertext[62]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_0_n3), .B(MCInst_MC3_v3_0[3]), .ZN(
        Red_SignaltoCheck[96]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_1_n3), .B(Red_MCInst_MC3_v3_1[2]), 
        .ZN(Red_SignaltoCheck[97]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_2_n3), .B(Red_MCInst_MC3_v3_1[2]), 
        .ZN(Red_SignaltoCheck[98]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_2_U1 ( .A(Red_MCInst_MC3_v3_3[2]), 
        .B(MCInst_MC3_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_0_n3), .B(MCInst_MC2_v3_0[3]), .ZN(
        Red_SignaltoCheck[99]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_1_n3), .B(Red_MCInst_MC2_v3_1[2]), 
        .ZN(Red_SignaltoCheck[100]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_2_n3), .B(Red_MCInst_MC2_v3_1[2]), 
        .ZN(Red_SignaltoCheck[101]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_2_U1 ( .A(Red_MCInst_MC2_v3_3[2]), 
        .B(MCInst_MC2_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_0_n3), .B(MCInst_MC1_v3_0[3]), .ZN(
        Red_SignaltoCheck[102]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_1_n3), .B(Red_MCInst_MC1_v3_1[2]), 
        .ZN(Red_SignaltoCheck[103]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_2_n3), .B(Red_MCInst_MC1_v3_1[2]), 
        .ZN(Red_SignaltoCheck[104]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_2_U1 ( .A(Red_MCInst_MC1_v3_3[2]), 
        .B(MCInst_MC1_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_0_n3), .B(MCInst_MC0_v3_0[3]), .ZN(
        Red_SignaltoCheck[105]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_1_n3), .B(Red_MCInst_MC0_v3_1[2]), 
        .ZN(Red_SignaltoCheck[106]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_2_n3), .B(Red_MCInst_MC0_v3_1[2]), 
        .ZN(Red_SignaltoCheck[107]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_2_U1 ( .A(Red_MCInst_MC0_v3_3[2]), 
        .B(MCInst_MC0_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_0_n3), .B(MCInst_MC3_v2_0[3]), .ZN(
        Red_SignaltoCheck[108]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U1 ( .A(ShiftRowsOutput[16]), 
        .B(MCInst_MC3_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_1_n3), .B(Red_MCInst_MC3_v2_2[1]), 
        .ZN(Red_SignaltoCheck[109]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_1_U1 ( .A(ShiftRowsOutput[16]), 
        .B(MCInst_MC3_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_2_n3), .B(Red_MCInst_MC3_v2_2[1]), 
        .ZN(Red_SignaltoCheck[110]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_2_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_0_n3), .B(MCInst_MC2_v2_0[3]), .ZN(
        Red_SignaltoCheck[111]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U1 ( .A(ShiftRowsOutput[20]), 
        .B(MCInst_MC2_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_1_n3), .B(Red_MCInst_MC2_v2_2[1]), 
        .ZN(Red_SignaltoCheck[112]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_1_U1 ( .A(ShiftRowsOutput[20]), 
        .B(MCInst_MC2_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_2_n3), .B(Red_MCInst_MC2_v2_2[1]), 
        .ZN(Red_SignaltoCheck[113]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_2_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_0_n3), .B(MCInst_MC1_v2_0[3]), .ZN(
        Red_SignaltoCheck[114]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U1 ( .A(ShiftRowsOutput[24]), 
        .B(MCInst_MC1_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_1_n3), .B(Red_MCInst_MC1_v2_2[1]), 
        .ZN(Red_SignaltoCheck[115]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_1_U1 ( .A(ShiftRowsOutput[24]), 
        .B(MCInst_MC1_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_2_n3), .B(Red_MCInst_MC1_v2_2[1]), 
        .ZN(Red_SignaltoCheck[116]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_2_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_0_n3), .B(MCInst_MC0_v2_0[3]), .ZN(
        Red_SignaltoCheck[117]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U1 ( .A(ShiftRowsOutput[28]), 
        .B(MCInst_MC0_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_1_n3), .B(Red_MCInst_MC0_v2_2[1]), 
        .ZN(Red_SignaltoCheck[118]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_1_U1 ( .A(ShiftRowsOutput[28]), 
        .B(MCInst_MC0_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_2_n3), .B(Red_MCInst_MC0_v2_2[1]), 
        .ZN(Red_SignaltoCheck[119]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_2_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_0_n3), .B(MCInst_MC3_v1_3[3]), .ZN(
        Red_SignaltoCheck[120]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_1_n3), .B(Red_MCInst_MC3_v1_1[2]), 
        .ZN(Red_SignaltoCheck[121]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_2_n3), .B(Red_MCInst_MC3_v1_1[2]), 
        .ZN(Red_SignaltoCheck[122]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_2_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        MCInst_MC3_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_0_n3), .B(MCInst_MC2_v1_3[3]), .ZN(
        Red_SignaltoCheck[123]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_1_n3), .B(Red_MCInst_MC2_v1_1[2]), 
        .ZN(Red_SignaltoCheck[124]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_2_n3), .B(Red_MCInst_MC2_v1_1[2]), 
        .ZN(Red_SignaltoCheck[125]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_2_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        MCInst_MC2_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_0_n3), .B(MCInst_MC1_v1_3[3]), .ZN(
        Red_SignaltoCheck[126]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_1_n3), .B(Red_MCInst_MC1_v1_1[2]), 
        .ZN(Red_SignaltoCheck[127]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_2_n3), .B(Red_MCInst_MC1_v1_1[2]), 
        .ZN(Red_SignaltoCheck[128]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_2_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        MCInst_MC1_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_0_n3), .B(MCInst_MC0_v1_3[3]), .ZN(
        Red_SignaltoCheck[129]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_1_n3), .B(Red_MCInst_MC0_v1_1[2]), 
        .ZN(Red_SignaltoCheck[130]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_2_n3), .B(Red_MCInst_MC0_v1_1[2]), 
        .ZN(Red_SignaltoCheck[131]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_2_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        MCInst_MC0_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_0_n3), .B(MCInst_MC3_v0_3[3]), .ZN(
        Red_SignaltoCheck[132]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), 
        .B(Red_MCInst_MC3_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_1_n3), .B(Red_MCInst_MC3_v0_1[0]), 
        .ZN(Red_SignaltoCheck[133]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), 
        .B(Red_MCInst_MC3_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_2_n3), .B(Red_MCInst_MC3_v0_1[0]), 
        .ZN(Red_SignaltoCheck[134]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), 
        .B(MCInst_MC3_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_0_n3), .B(MCInst_MC2_v0_3[3]), .ZN(
        Red_SignaltoCheck[135]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), 
        .B(Red_MCInst_MC2_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_1_n3), .B(Red_MCInst_MC2_v0_1[0]), 
        .ZN(Red_SignaltoCheck[136]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), 
        .B(Red_MCInst_MC2_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_2_n3), .B(Red_MCInst_MC2_v0_1[0]), 
        .ZN(Red_SignaltoCheck[137]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), 
        .B(MCInst_MC2_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_0_n3), .B(MCInst_MC1_v0_3[3]), .ZN(
        Red_SignaltoCheck[138]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), 
        .B(Red_MCInst_MC1_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_1_n3), .B(Red_MCInst_MC1_v0_1[0]), 
        .ZN(Red_SignaltoCheck[139]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), 
        .B(Red_MCInst_MC1_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_2_n3), .B(Red_MCInst_MC1_v0_1[0]), 
        .ZN(Red_SignaltoCheck[140]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), 
        .B(MCInst_MC1_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_0_n3), .B(MCInst_MC0_v0_3[3]), .ZN(
        Red_SignaltoCheck[141]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), 
        .B(Red_MCInst_MC0_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_1_n3), .B(Red_MCInst_MC0_v0_1[0]), 
        .ZN(Red_SignaltoCheck[142]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), 
        .B(Red_MCInst_MC0_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_2_n3), .B(Red_MCInst_MC0_v0_1[0]), 
        .ZN(Red_SignaltoCheck[143]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), 
        .B(MCInst_MC0_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_2_n3) );
  NOR2_X1 Check1_CheckInst_0_U95 ( .A1(Check1_CheckInst_0_n94), .A2(
        Check1_CheckInst_0_n93), .ZN(Error[0]) );
  NAND2_X1 Check1_CheckInst_0_U94 ( .A1(Check1_CheckInst_0_n92), .A2(
        Check1_CheckInst_0_n91), .ZN(Check1_CheckInst_0_n93) );
  NOR2_X1 Check1_CheckInst_0_U93 ( .A1(Check1_CheckInst_0_n90), .A2(
        Check1_CheckInst_0_n89), .ZN(Check1_CheckInst_0_n91) );
  NAND2_X1 Check1_CheckInst_0_U92 ( .A1(Check1_CheckInst_0_n88), .A2(
        Check1_CheckInst_0_n87), .ZN(Check1_CheckInst_0_n89) );
  NOR2_X1 Check1_CheckInst_0_U91 ( .A1(Check1_CheckInst_0_n86), .A2(
        Check1_CheckInst_0_n85), .ZN(Check1_CheckInst_0_n87) );
  NAND2_X1 Check1_CheckInst_0_U90 ( .A1(Check1_CheckInst_0_n84), .A2(
        Check1_CheckInst_0_n83), .ZN(Check1_CheckInst_0_n85) );
  NOR2_X1 Check1_CheckInst_0_U89 ( .A1(Check1_CheckInst_0_n82), .A2(
        Check1_CheckInst_0_n81), .ZN(Check1_CheckInst_0_n83) );
  XOR2_X1 Check1_CheckInst_0_U88 ( .A(Red_AddRoundKeyOutput[21]), .B(
        Red_SignaltoCheck[21]), .Z(Check1_CheckInst_0_n81) );
  XOR2_X1 Check1_CheckInst_0_U87 ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[15]), .Z(Check1_CheckInst_0_n82) );
  XNOR2_X1 Check1_CheckInst_0_U86 ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[9]), .ZN(Check1_CheckInst_0_n84) );
  NAND2_X1 Check1_CheckInst_0_U85 ( .A1(Check1_CheckInst_0_n80), .A2(
        Check1_CheckInst_0_n79), .ZN(Check1_CheckInst_0_n86) );
  NOR2_X1 Check1_CheckInst_0_U84 ( .A1(Check1_CheckInst_0_n78), .A2(
        Check1_CheckInst_0_n77), .ZN(Check1_CheckInst_0_n79) );
  NAND2_X1 Check1_CheckInst_0_U83 ( .A1(Check1_CheckInst_0_n76), .A2(
        Check1_CheckInst_0_n75), .ZN(Check1_CheckInst_0_n77) );
  NOR2_X1 Check1_CheckInst_0_U82 ( .A1(Check1_CheckInst_0_n74), .A2(
        Check1_CheckInst_0_n73), .ZN(Check1_CheckInst_0_n75) );
  XOR2_X1 Check1_CheckInst_0_U81 ( .A(Red_AddRoundKeyOutput[24]), .B(
        Red_SignaltoCheck[24]), .Z(Check1_CheckInst_0_n73) );
  XOR2_X1 Check1_CheckInst_0_U80 ( .A(Red_AddRoundKeyOutput[27]), .B(
        Red_SignaltoCheck[27]), .Z(Check1_CheckInst_0_n74) );
  XNOR2_X1 Check1_CheckInst_0_U79 ( .A(Red_AddRoundKeyOutput[30]), .B(
        Red_SignaltoCheck[30]), .ZN(Check1_CheckInst_0_n76) );
  NAND2_X1 Check1_CheckInst_0_U78 ( .A1(Check1_CheckInst_0_n72), .A2(
        Check1_CheckInst_0_n71), .ZN(Check1_CheckInst_0_n78) );
  NOR2_X1 Check1_CheckInst_0_U77 ( .A1(Check1_CheckInst_0_n70), .A2(
        Check1_CheckInst_0_n69), .ZN(Check1_CheckInst_0_n71) );
  NAND2_X1 Check1_CheckInst_0_U76 ( .A1(Check1_CheckInst_0_n68), .A2(
        Check1_CheckInst_0_n67), .ZN(Check1_CheckInst_0_n69) );
  NOR2_X1 Check1_CheckInst_0_U75 ( .A1(Check1_CheckInst_0_n66), .A2(
        Check1_CheckInst_0_n65), .ZN(Check1_CheckInst_0_n67) );
  XOR2_X1 Check1_CheckInst_0_U74 ( .A(Red_ShiftRowsOutput[12]), .B(
        Red_SignaltoCheck[108]), .Z(Check1_CheckInst_0_n65) );
  XOR2_X1 Check1_CheckInst_0_U73 ( .A(Red_ShiftRowsOutput[24]), .B(
        Red_SignaltoCheck[120]), .Z(Check1_CheckInst_0_n66) );
  XNOR2_X1 Check1_CheckInst_0_U72 ( .A(Red_ShiftRowsOutput[9]), .B(
        Red_SignaltoCheck[105]), .ZN(Check1_CheckInst_0_n68) );
  NAND2_X1 Check1_CheckInst_0_U71 ( .A1(Check1_CheckInst_0_n64), .A2(
        Check1_CheckInst_0_n63), .ZN(Check1_CheckInst_0_n70) );
  NOR2_X1 Check1_CheckInst_0_U70 ( .A1(Check1_CheckInst_0_n62), .A2(
        Check1_CheckInst_0_n61), .ZN(Check1_CheckInst_0_n63) );
  XOR2_X1 Check1_CheckInst_0_U69 ( .A(Red_ShiftRowsOutput[18]), .B(
        Red_SignaltoCheck[114]), .Z(Check1_CheckInst_0_n61) );
  XOR2_X1 Check1_CheckInst_0_U68 ( .A(Red_ShiftRowsOutput[21]), .B(
        Red_SignaltoCheck[117]), .Z(Check1_CheckInst_0_n62) );
  NOR2_X1 Check1_CheckInst_0_U67 ( .A1(Check1_CheckInst_0_n60), .A2(
        Check1_CheckInst_0_n59), .ZN(Check1_CheckInst_0_n64) );
  XOR2_X1 Check1_CheckInst_0_U66 ( .A(Red_ShiftRowsOutput[33]), .B(
        Red_SignaltoCheck[129]), .Z(Check1_CheckInst_0_n59) );
  XOR2_X1 Check1_CheckInst_0_U65 ( .A(Red_ShiftRowsOutput[27]), .B(
        Red_SignaltoCheck[123]), .Z(Check1_CheckInst_0_n60) );
  XNOR2_X1 Check1_CheckInst_0_U64 ( .A(Red_SignaltoCheck[111]), .B(
        Red_ShiftRowsOutput[15]), .ZN(Check1_CheckInst_0_n72) );
  XNOR2_X1 Check1_CheckInst_0_U63 ( .A(Red_SignaltoCheck[18]), .B(
        Red_AddRoundKeyOutput[18]), .ZN(Check1_CheckInst_0_n80) );
  XNOR2_X1 Check1_CheckInst_0_U62 ( .A(Red_SignaltoCheck[6]), .B(
        Red_AddRoundKeyOutput[6]), .ZN(Check1_CheckInst_0_n88) );
  NAND2_X1 Check1_CheckInst_0_U61 ( .A1(Check1_CheckInst_0_n58), .A2(
        Check1_CheckInst_0_n57), .ZN(Check1_CheckInst_0_n90) );
  NOR2_X1 Check1_CheckInst_0_U60 ( .A1(Check1_CheckInst_0_n56), .A2(
        Check1_CheckInst_0_n55), .ZN(Check1_CheckInst_0_n57) );
  NAND2_X1 Check1_CheckInst_0_U59 ( .A1(Check1_CheckInst_0_n54), .A2(
        Check1_CheckInst_0_n53), .ZN(Check1_CheckInst_0_n55) );
  NOR2_X1 Check1_CheckInst_0_U58 ( .A1(Check1_CheckInst_0_n52), .A2(
        Check1_CheckInst_0_n51), .ZN(Check1_CheckInst_0_n53) );
  XOR2_X1 Check1_CheckInst_0_U57 ( .A(Red_AddRoundKeyOutput[36]), .B(
        Red_SignaltoCheck[36]), .Z(Check1_CheckInst_0_n51) );
  XOR2_X1 Check1_CheckInst_0_U56 ( .A(Red_MC_output[0]), .B(
        Red_SignaltoCheck[48]), .Z(Check1_CheckInst_0_n52) );
  XNOR2_X1 Check1_CheckInst_0_U55 ( .A(Red_AddRoundKeyOutput[33]), .B(
        Red_SignaltoCheck[33]), .ZN(Check1_CheckInst_0_n54) );
  NAND2_X1 Check1_CheckInst_0_U54 ( .A1(Check1_CheckInst_0_n50), .A2(
        Check1_CheckInst_0_n49), .ZN(Check1_CheckInst_0_n56) );
  NOR2_X1 Check1_CheckInst_0_U53 ( .A1(Check1_CheckInst_0_n48), .A2(
        Check1_CheckInst_0_n47), .ZN(Check1_CheckInst_0_n49) );
  NAND2_X1 Check1_CheckInst_0_U52 ( .A1(Check1_CheckInst_0_n46), .A2(
        Check1_CheckInst_0_n45), .ZN(Check1_CheckInst_0_n47) );
  NOR2_X1 Check1_CheckInst_0_U51 ( .A1(Check1_CheckInst_0_n44), .A2(
        Check1_CheckInst_0_n43), .ZN(Check1_CheckInst_0_n45) );
  XOR2_X1 Check1_CheckInst_0_U50 ( .A(Red_MC_output[9]), .B(
        Red_SignaltoCheck[57]), .Z(Check1_CheckInst_0_n43) );
  XOR2_X1 Check1_CheckInst_0_U49 ( .A(Red_MC_output[3]), .B(
        Red_SignaltoCheck[51]), .Z(Check1_CheckInst_0_n44) );
  XNOR2_X1 Check1_CheckInst_0_U48 ( .A(Red_AddRoundKeyOutput[45]), .B(
        Red_SignaltoCheck[45]), .ZN(Check1_CheckInst_0_n46) );
  NAND2_X1 Check1_CheckInst_0_U47 ( .A1(Check1_CheckInst_0_n42), .A2(
        Check1_CheckInst_0_n41), .ZN(Check1_CheckInst_0_n48) );
  NOR2_X1 Check1_CheckInst_0_U46 ( .A1(Check1_CheckInst_0_n40), .A2(
        Check1_CheckInst_0_n39), .ZN(Check1_CheckInst_0_n41) );
  NAND2_X1 Check1_CheckInst_0_U45 ( .A1(Check1_CheckInst_0_n38), .A2(
        Check1_CheckInst_0_n37), .ZN(Check1_CheckInst_0_n39) );
  NOR2_X1 Check1_CheckInst_0_U44 ( .A1(Check1_CheckInst_0_n36), .A2(
        Check1_CheckInst_0_n35), .ZN(Check1_CheckInst_0_n37) );
  XOR2_X1 Check1_CheckInst_0_U43 ( .A(Red_MC_output[12]), .B(
        Red_SignaltoCheck[60]), .Z(Check1_CheckInst_0_n35) );
  XOR2_X1 Check1_CheckInst_0_U42 ( .A(Red_MC_output[15]), .B(
        Red_SignaltoCheck[63]), .Z(Check1_CheckInst_0_n36) );
  XNOR2_X1 Check1_CheckInst_0_U41 ( .A(Red_MC_output[18]), .B(
        Red_SignaltoCheck[66]), .ZN(Check1_CheckInst_0_n38) );
  NAND2_X1 Check1_CheckInst_0_U40 ( .A1(Check1_CheckInst_0_n34), .A2(
        Check1_CheckInst_0_n33), .ZN(Check1_CheckInst_0_n40) );
  NOR2_X1 Check1_CheckInst_0_U39 ( .A1(Check1_CheckInst_0_n32), .A2(
        Check1_CheckInst_0_n31), .ZN(Check1_CheckInst_0_n33) );
  XOR2_X1 Check1_CheckInst_0_U38 ( .A(Red_ShiftRowsOutput[45]), .B(
        Red_SignaltoCheck[141]), .Z(Check1_CheckInst_0_n31) );
  XOR2_X1 Check1_CheckInst_0_U37 ( .A(Red_SignaltoCheck[3]), .B(
        Red_AddRoundKeyOutput[3]), .Z(Check1_CheckInst_0_n32) );
  NOR2_X1 Check1_CheckInst_0_U36 ( .A1(Check1_CheckInst_0_n30), .A2(
        Check1_CheckInst_0_n29), .ZN(Check1_CheckInst_0_n34) );
  XOR2_X1 Check1_CheckInst_0_U35 ( .A(Red_AddRoundKeyOutput[0]), .B(
        Red_SignaltoCheck[0]), .Z(Check1_CheckInst_0_n29) );
  XOR2_X1 Check1_CheckInst_0_U34 ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[12]), .Z(Check1_CheckInst_0_n30) );
  XNOR2_X1 Check1_CheckInst_0_U33 ( .A(Red_SignaltoCheck[54]), .B(
        Red_MC_output[6]), .ZN(Check1_CheckInst_0_n42) );
  XNOR2_X1 Check1_CheckInst_0_U32 ( .A(Red_SignaltoCheck[42]), .B(
        Red_AddRoundKeyOutput[42]), .ZN(Check1_CheckInst_0_n50) );
  XNOR2_X1 Check1_CheckInst_0_U31 ( .A(Red_SignaltoCheck[39]), .B(
        Red_AddRoundKeyOutput[39]), .ZN(Check1_CheckInst_0_n58) );
  NOR2_X1 Check1_CheckInst_0_U30 ( .A1(Check1_CheckInst_0_n28), .A2(
        Check1_CheckInst_0_n27), .ZN(Check1_CheckInst_0_n92) );
  NAND2_X1 Check1_CheckInst_0_U29 ( .A1(Check1_CheckInst_0_n26), .A2(
        Check1_CheckInst_0_n25), .ZN(Check1_CheckInst_0_n27) );
  NOR2_X1 Check1_CheckInst_0_U28 ( .A1(Check1_CheckInst_0_n24), .A2(
        Check1_CheckInst_0_n23), .ZN(Check1_CheckInst_0_n25) );
  NAND2_X1 Check1_CheckInst_0_U27 ( .A1(Check1_CheckInst_0_n22), .A2(
        Check1_CheckInst_0_n21), .ZN(Check1_CheckInst_0_n23) );
  XNOR2_X1 Check1_CheckInst_0_U26 ( .A(Red_ShiftRowsOutput[0]), .B(
        Red_SignaltoCheck[96]), .ZN(Check1_CheckInst_0_n21) );
  XNOR2_X1 Check1_CheckInst_0_U25 ( .A(Red_ShiftRowsOutput[3]), .B(
        Red_SignaltoCheck[99]), .ZN(Check1_CheckInst_0_n22) );
  NAND2_X1 Check1_CheckInst_0_U24 ( .A1(Check1_CheckInst_0_n20), .A2(
        Check1_CheckInst_0_n19), .ZN(Check1_CheckInst_0_n24) );
  XNOR2_X1 Check1_CheckInst_0_U23 ( .A(Red_MC_output[42]), .B(
        Red_SignaltoCheck[90]), .ZN(Check1_CheckInst_0_n19) );
  XNOR2_X1 Check1_CheckInst_0_U22 ( .A(Red_ShiftRowsOutput[6]), .B(
        Red_SignaltoCheck[102]), .ZN(Check1_CheckInst_0_n20) );
  NOR2_X1 Check1_CheckInst_0_U21 ( .A1(Check1_CheckInst_0_n18), .A2(
        Check1_CheckInst_0_n17), .ZN(Check1_CheckInst_0_n26) );
  XOR2_X1 Check1_CheckInst_0_U20 ( .A(Red_MC_output[45]), .B(
        Red_SignaltoCheck[93]), .Z(Check1_CheckInst_0_n17) );
  XOR2_X1 Check1_CheckInst_0_U19 ( .A(Red_MC_output[39]), .B(
        Red_SignaltoCheck[87]), .Z(Check1_CheckInst_0_n18) );
  NAND2_X1 Check1_CheckInst_0_U18 ( .A1(Check1_CheckInst_0_n16), .A2(
        Check1_CheckInst_0_n15), .ZN(Check1_CheckInst_0_n28) );
  XNOR2_X1 Check1_CheckInst_0_U17 ( .A(Red_MC_output[30]), .B(
        Red_SignaltoCheck[78]), .ZN(Check1_CheckInst_0_n15) );
  XNOR2_X1 Check1_CheckInst_0_U16 ( .A(Red_MC_output[33]), .B(
        Red_SignaltoCheck[81]), .ZN(Check1_CheckInst_0_n16) );
  NAND2_X1 Check1_CheckInst_0_U15 ( .A1(Check1_CheckInst_0_n14), .A2(
        Check1_CheckInst_0_n13), .ZN(Check1_CheckInst_0_n94) );
  NOR2_X1 Check1_CheckInst_0_U14 ( .A1(Check1_CheckInst_0_n12), .A2(
        Check1_CheckInst_0_n11), .ZN(Check1_CheckInst_0_n13) );
  NAND2_X1 Check1_CheckInst_0_U13 ( .A1(Check1_CheckInst_0_n10), .A2(
        Check1_CheckInst_0_n9), .ZN(Check1_CheckInst_0_n11) );
  NOR2_X1 Check1_CheckInst_0_U12 ( .A1(Check1_CheckInst_0_n8), .A2(
        Check1_CheckInst_0_n7), .ZN(Check1_CheckInst_0_n9) );
  XOR2_X1 Check1_CheckInst_0_U11 ( .A(Red_MC_output[24]), .B(
        Red_SignaltoCheck[72]), .Z(Check1_CheckInst_0_n7) );
  XOR2_X1 Check1_CheckInst_0_U10 ( .A(Red_MC_output[36]), .B(
        Red_SignaltoCheck[84]), .Z(Check1_CheckInst_0_n8) );
  NOR2_X1 Check1_CheckInst_0_U9 ( .A1(Check1_CheckInst_0_n6), .A2(
        Check1_CheckInst_0_n5), .ZN(Check1_CheckInst_0_n10) );
  XOR2_X1 Check1_CheckInst_0_U8 ( .A(Red_MC_output[27]), .B(
        Red_SignaltoCheck[75]), .Z(Check1_CheckInst_0_n5) );
  XOR2_X1 Check1_CheckInst_0_U7 ( .A(Red_MC_output[21]), .B(
        Red_SignaltoCheck[69]), .Z(Check1_CheckInst_0_n6) );
  NAND2_X1 Check1_CheckInst_0_U6 ( .A1(Check1_CheckInst_0_n4), .A2(
        Check1_CheckInst_0_n3), .ZN(Check1_CheckInst_0_n12) );
  XNOR2_X1 Check1_CheckInst_0_U5 ( .A(Red_ShiftRowsOutput[36]), .B(
        Red_SignaltoCheck[132]), .ZN(Check1_CheckInst_0_n3) );
  XNOR2_X1 Check1_CheckInst_0_U4 ( .A(Red_ShiftRowsOutput[39]), .B(
        Red_SignaltoCheck[135]), .ZN(Check1_CheckInst_0_n4) );
  NOR2_X1 Check1_CheckInst_0_U3 ( .A1(Check1_CheckInst_0_n2), .A2(
        Check1_CheckInst_0_n1), .ZN(Check1_CheckInst_0_n14) );
  XOR2_X1 Check1_CheckInst_0_U2 ( .A(Red_ShiftRowsOutput[30]), .B(
        Red_SignaltoCheck[126]), .Z(Check1_CheckInst_0_n1) );
  XOR2_X1 Check1_CheckInst_0_U1 ( .A(Red_ShiftRowsOutput[42]), .B(
        Red_SignaltoCheck[138]), .Z(Check1_CheckInst_0_n2) );
  NOR2_X1 Check1_CheckInst_1_U95 ( .A1(Check1_CheckInst_1_n96), .A2(
        Check1_CheckInst_1_n95), .ZN(Error[1]) );
  NAND2_X1 Check1_CheckInst_1_U94 ( .A1(Check1_CheckInst_1_n94), .A2(
        Check1_CheckInst_1_n93), .ZN(Check1_CheckInst_1_n95) );
  NOR2_X1 Check1_CheckInst_1_U93 ( .A1(Check1_CheckInst_1_n92), .A2(
        Check1_CheckInst_1_n91), .ZN(Check1_CheckInst_1_n93) );
  NAND2_X1 Check1_CheckInst_1_U92 ( .A1(Check1_CheckInst_1_n90), .A2(
        Check1_CheckInst_1_n89), .ZN(Check1_CheckInst_1_n91) );
  NOR2_X1 Check1_CheckInst_1_U91 ( .A1(Check1_CheckInst_1_n88), .A2(
        Check1_CheckInst_1_n87), .ZN(Check1_CheckInst_1_n89) );
  NAND2_X1 Check1_CheckInst_1_U90 ( .A1(Check1_CheckInst_1_n86), .A2(
        Check1_CheckInst_1_n85), .ZN(Check1_CheckInst_1_n87) );
  NOR2_X1 Check1_CheckInst_1_U89 ( .A1(Check1_CheckInst_1_n84), .A2(
        Check1_CheckInst_1_n83), .ZN(Check1_CheckInst_1_n85) );
  XOR2_X1 Check1_CheckInst_1_U88 ( .A(Red_AddRoundKeyOutput[22]), .B(
        Red_SignaltoCheck[22]), .Z(Check1_CheckInst_1_n83) );
  XOR2_X1 Check1_CheckInst_1_U87 ( .A(Red_AddRoundKeyOutput[16]), .B(
        Red_SignaltoCheck[16]), .Z(Check1_CheckInst_1_n84) );
  XNOR2_X1 Check1_CheckInst_1_U86 ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[10]), .ZN(Check1_CheckInst_1_n86) );
  NAND2_X1 Check1_CheckInst_1_U85 ( .A1(Check1_CheckInst_1_n82), .A2(
        Check1_CheckInst_1_n81), .ZN(Check1_CheckInst_1_n88) );
  NOR2_X1 Check1_CheckInst_1_U84 ( .A1(Check1_CheckInst_1_n80), .A2(
        Check1_CheckInst_1_n79), .ZN(Check1_CheckInst_1_n81) );
  NAND2_X1 Check1_CheckInst_1_U83 ( .A1(Check1_CheckInst_1_n78), .A2(
        Check1_CheckInst_1_n77), .ZN(Check1_CheckInst_1_n79) );
  NOR2_X1 Check1_CheckInst_1_U82 ( .A1(Check1_CheckInst_1_n76), .A2(
        Check1_CheckInst_1_n75), .ZN(Check1_CheckInst_1_n77) );
  XOR2_X1 Check1_CheckInst_1_U81 ( .A(Red_AddRoundKeyOutput[25]), .B(
        Red_SignaltoCheck[25]), .Z(Check1_CheckInst_1_n75) );
  XOR2_X1 Check1_CheckInst_1_U80 ( .A(Red_AddRoundKeyOutput[28]), .B(
        Red_SignaltoCheck[28]), .Z(Check1_CheckInst_1_n76) );
  XNOR2_X1 Check1_CheckInst_1_U79 ( .A(Red_AddRoundKeyOutput[31]), .B(
        Red_SignaltoCheck[31]), .ZN(Check1_CheckInst_1_n78) );
  NAND2_X1 Check1_CheckInst_1_U78 ( .A1(Check1_CheckInst_1_n74), .A2(
        Check1_CheckInst_1_n73), .ZN(Check1_CheckInst_1_n80) );
  NOR2_X1 Check1_CheckInst_1_U77 ( .A1(Check1_CheckInst_1_n72), .A2(
        Check1_CheckInst_1_n71), .ZN(Check1_CheckInst_1_n73) );
  NAND2_X1 Check1_CheckInst_1_U76 ( .A1(Check1_CheckInst_1_n70), .A2(
        Check1_CheckInst_1_n69), .ZN(Check1_CheckInst_1_n71) );
  NOR2_X1 Check1_CheckInst_1_U75 ( .A1(Check1_CheckInst_1_n68), .A2(
        Check1_CheckInst_1_n67), .ZN(Check1_CheckInst_1_n69) );
  XOR2_X1 Check1_CheckInst_1_U74 ( .A(Red_ShiftRowsOutput[13]), .B(
        Red_SignaltoCheck[109]), .Z(Check1_CheckInst_1_n67) );
  XOR2_X1 Check1_CheckInst_1_U73 ( .A(Red_ShiftRowsOutput[25]), .B(
        Red_SignaltoCheck[121]), .Z(Check1_CheckInst_1_n68) );
  XNOR2_X1 Check1_CheckInst_1_U72 ( .A(Red_ShiftRowsOutput[10]), .B(
        Red_SignaltoCheck[106]), .ZN(Check1_CheckInst_1_n70) );
  NAND2_X1 Check1_CheckInst_1_U71 ( .A1(Check1_CheckInst_1_n66), .A2(
        Check1_CheckInst_1_n65), .ZN(Check1_CheckInst_1_n72) );
  NOR2_X1 Check1_CheckInst_1_U70 ( .A1(Check1_CheckInst_1_n64), .A2(
        Check1_CheckInst_1_n63), .ZN(Check1_CheckInst_1_n65) );
  XOR2_X1 Check1_CheckInst_1_U69 ( .A(Red_ShiftRowsOutput[19]), .B(
        Red_SignaltoCheck[115]), .Z(Check1_CheckInst_1_n63) );
  XOR2_X1 Check1_CheckInst_1_U68 ( .A(Red_ShiftRowsOutput[22]), .B(
        Red_SignaltoCheck[118]), .Z(Check1_CheckInst_1_n64) );
  NOR2_X1 Check1_CheckInst_1_U67 ( .A1(Check1_CheckInst_1_n62), .A2(
        Check1_CheckInst_1_n61), .ZN(Check1_CheckInst_1_n66) );
  XOR2_X1 Check1_CheckInst_1_U66 ( .A(Red_ShiftRowsOutput[34]), .B(
        Red_SignaltoCheck[130]), .Z(Check1_CheckInst_1_n61) );
  XOR2_X1 Check1_CheckInst_1_U65 ( .A(Red_ShiftRowsOutput[28]), .B(
        Red_SignaltoCheck[124]), .Z(Check1_CheckInst_1_n62) );
  XNOR2_X1 Check1_CheckInst_1_U64 ( .A(Red_SignaltoCheck[112]), .B(
        Red_ShiftRowsOutput[16]), .ZN(Check1_CheckInst_1_n74) );
  XNOR2_X1 Check1_CheckInst_1_U63 ( .A(Red_SignaltoCheck[19]), .B(
        Red_AddRoundKeyOutput[19]), .ZN(Check1_CheckInst_1_n82) );
  XNOR2_X1 Check1_CheckInst_1_U62 ( .A(Red_SignaltoCheck[7]), .B(
        Red_AddRoundKeyOutput[7]), .ZN(Check1_CheckInst_1_n90) );
  NAND2_X1 Check1_CheckInst_1_U61 ( .A1(Check1_CheckInst_1_n60), .A2(
        Check1_CheckInst_1_n59), .ZN(Check1_CheckInst_1_n92) );
  NOR2_X1 Check1_CheckInst_1_U60 ( .A1(Check1_CheckInst_1_n58), .A2(
        Check1_CheckInst_1_n57), .ZN(Check1_CheckInst_1_n59) );
  NAND2_X1 Check1_CheckInst_1_U59 ( .A1(Check1_CheckInst_1_n56), .A2(
        Check1_CheckInst_1_n55), .ZN(Check1_CheckInst_1_n57) );
  NOR2_X1 Check1_CheckInst_1_U58 ( .A1(Check1_CheckInst_1_n54), .A2(
        Check1_CheckInst_1_n53), .ZN(Check1_CheckInst_1_n55) );
  XOR2_X1 Check1_CheckInst_1_U57 ( .A(Red_AddRoundKeyOutput[37]), .B(
        Red_SignaltoCheck[37]), .Z(Check1_CheckInst_1_n53) );
  XOR2_X1 Check1_CheckInst_1_U56 ( .A(Red_MC_output[1]), .B(
        Red_SignaltoCheck[49]), .Z(Check1_CheckInst_1_n54) );
  XNOR2_X1 Check1_CheckInst_1_U55 ( .A(Red_AddRoundKeyOutput[34]), .B(
        Red_SignaltoCheck[34]), .ZN(Check1_CheckInst_1_n56) );
  NAND2_X1 Check1_CheckInst_1_U54 ( .A1(Check1_CheckInst_1_n52), .A2(
        Check1_CheckInst_1_n51), .ZN(Check1_CheckInst_1_n58) );
  NOR2_X1 Check1_CheckInst_1_U53 ( .A1(Check1_CheckInst_1_n50), .A2(
        Check1_CheckInst_1_n49), .ZN(Check1_CheckInst_1_n51) );
  NAND2_X1 Check1_CheckInst_1_U52 ( .A1(Check1_CheckInst_1_n48), .A2(
        Check1_CheckInst_1_n47), .ZN(Check1_CheckInst_1_n49) );
  NOR2_X1 Check1_CheckInst_1_U51 ( .A1(Check1_CheckInst_1_n46), .A2(
        Check1_CheckInst_1_n45), .ZN(Check1_CheckInst_1_n47) );
  XOR2_X1 Check1_CheckInst_1_U50 ( .A(Red_MC_output[10]), .B(
        Red_SignaltoCheck[58]), .Z(Check1_CheckInst_1_n45) );
  XOR2_X1 Check1_CheckInst_1_U49 ( .A(Red_MC_output[4]), .B(
        Red_SignaltoCheck[52]), .Z(Check1_CheckInst_1_n46) );
  XNOR2_X1 Check1_CheckInst_1_U48 ( .A(Red_AddRoundKeyOutput[46]), .B(
        Red_SignaltoCheck[46]), .ZN(Check1_CheckInst_1_n48) );
  NAND2_X1 Check1_CheckInst_1_U47 ( .A1(Check1_CheckInst_1_n44), .A2(
        Check1_CheckInst_1_n43), .ZN(Check1_CheckInst_1_n50) );
  NOR2_X1 Check1_CheckInst_1_U46 ( .A1(Check1_CheckInst_1_n42), .A2(
        Check1_CheckInst_1_n41), .ZN(Check1_CheckInst_1_n43) );
  NAND2_X1 Check1_CheckInst_1_U45 ( .A1(Check1_CheckInst_1_n40), .A2(
        Check1_CheckInst_1_n39), .ZN(Check1_CheckInst_1_n41) );
  NOR2_X1 Check1_CheckInst_1_U44 ( .A1(Check1_CheckInst_1_n38), .A2(
        Check1_CheckInst_1_n37), .ZN(Check1_CheckInst_1_n39) );
  XOR2_X1 Check1_CheckInst_1_U43 ( .A(Red_MC_output[13]), .B(
        Red_SignaltoCheck[61]), .Z(Check1_CheckInst_1_n37) );
  XOR2_X1 Check1_CheckInst_1_U42 ( .A(Red_MC_output[16]), .B(
        Red_SignaltoCheck[64]), .Z(Check1_CheckInst_1_n38) );
  XNOR2_X1 Check1_CheckInst_1_U41 ( .A(Red_MC_output[19]), .B(
        Red_SignaltoCheck[67]), .ZN(Check1_CheckInst_1_n40) );
  NAND2_X1 Check1_CheckInst_1_U40 ( .A1(Check1_CheckInst_1_n36), .A2(
        Check1_CheckInst_1_n35), .ZN(Check1_CheckInst_1_n42) );
  NOR2_X1 Check1_CheckInst_1_U39 ( .A1(Check1_CheckInst_1_n34), .A2(
        Check1_CheckInst_1_n33), .ZN(Check1_CheckInst_1_n35) );
  XOR2_X1 Check1_CheckInst_1_U38 ( .A(Red_ShiftRowsOutput[46]), .B(
        Red_SignaltoCheck[142]), .Z(Check1_CheckInst_1_n33) );
  XOR2_X1 Check1_CheckInst_1_U37 ( .A(Red_SignaltoCheck[4]), .B(
        Red_AddRoundKeyOutput[4]), .Z(Check1_CheckInst_1_n34) );
  NOR2_X1 Check1_CheckInst_1_U36 ( .A1(Check1_CheckInst_1_n32), .A2(
        Check1_CheckInst_1_n31), .ZN(Check1_CheckInst_1_n36) );
  XOR2_X1 Check1_CheckInst_1_U35 ( .A(Red_AddRoundKeyOutput[1]), .B(
        Red_SignaltoCheck[1]), .Z(Check1_CheckInst_1_n31) );
  XOR2_X1 Check1_CheckInst_1_U34 ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[13]), .Z(Check1_CheckInst_1_n32) );
  XNOR2_X1 Check1_CheckInst_1_U33 ( .A(Red_SignaltoCheck[55]), .B(
        Red_MC_output[7]), .ZN(Check1_CheckInst_1_n44) );
  XNOR2_X1 Check1_CheckInst_1_U32 ( .A(Red_SignaltoCheck[43]), .B(
        Red_AddRoundKeyOutput[43]), .ZN(Check1_CheckInst_1_n52) );
  XNOR2_X1 Check1_CheckInst_1_U31 ( .A(Red_SignaltoCheck[40]), .B(
        Red_AddRoundKeyOutput[40]), .ZN(Check1_CheckInst_1_n60) );
  NOR2_X1 Check1_CheckInst_1_U30 ( .A1(Check1_CheckInst_1_n30), .A2(
        Check1_CheckInst_1_n29), .ZN(Check1_CheckInst_1_n94) );
  NAND2_X1 Check1_CheckInst_1_U29 ( .A1(Check1_CheckInst_1_n28), .A2(
        Check1_CheckInst_1_n27), .ZN(Check1_CheckInst_1_n29) );
  NOR2_X1 Check1_CheckInst_1_U28 ( .A1(Check1_CheckInst_1_n26), .A2(
        Check1_CheckInst_1_n25), .ZN(Check1_CheckInst_1_n27) );
  NAND2_X1 Check1_CheckInst_1_U27 ( .A1(Check1_CheckInst_1_n24), .A2(
        Check1_CheckInst_1_n23), .ZN(Check1_CheckInst_1_n25) );
  XNOR2_X1 Check1_CheckInst_1_U26 ( .A(Red_ShiftRowsOutput[1]), .B(
        Red_SignaltoCheck[97]), .ZN(Check1_CheckInst_1_n23) );
  XNOR2_X1 Check1_CheckInst_1_U25 ( .A(Red_ShiftRowsOutput[4]), .B(
        Red_SignaltoCheck[100]), .ZN(Check1_CheckInst_1_n24) );
  NAND2_X1 Check1_CheckInst_1_U24 ( .A1(Check1_CheckInst_1_n22), .A2(
        Check1_CheckInst_1_n21), .ZN(Check1_CheckInst_1_n26) );
  XNOR2_X1 Check1_CheckInst_1_U23 ( .A(Red_MC_output[43]), .B(
        Red_SignaltoCheck[91]), .ZN(Check1_CheckInst_1_n21) );
  XNOR2_X1 Check1_CheckInst_1_U22 ( .A(Red_ShiftRowsOutput[7]), .B(
        Red_SignaltoCheck[103]), .ZN(Check1_CheckInst_1_n22) );
  NOR2_X1 Check1_CheckInst_1_U21 ( .A1(Check1_CheckInst_1_n20), .A2(
        Check1_CheckInst_1_n19), .ZN(Check1_CheckInst_1_n28) );
  XOR2_X1 Check1_CheckInst_1_U20 ( .A(Red_MC_output[46]), .B(
        Red_SignaltoCheck[94]), .Z(Check1_CheckInst_1_n19) );
  XOR2_X1 Check1_CheckInst_1_U19 ( .A(Red_MC_output[40]), .B(
        Red_SignaltoCheck[88]), .Z(Check1_CheckInst_1_n20) );
  NAND2_X1 Check1_CheckInst_1_U18 ( .A1(Check1_CheckInst_1_n18), .A2(
        Check1_CheckInst_1_n17), .ZN(Check1_CheckInst_1_n30) );
  XNOR2_X1 Check1_CheckInst_1_U17 ( .A(Red_MC_output[31]), .B(
        Red_SignaltoCheck[79]), .ZN(Check1_CheckInst_1_n17) );
  XNOR2_X1 Check1_CheckInst_1_U16 ( .A(Red_MC_output[34]), .B(
        Red_SignaltoCheck[82]), .ZN(Check1_CheckInst_1_n18) );
  NAND2_X1 Check1_CheckInst_1_U15 ( .A1(Check1_CheckInst_1_n16), .A2(
        Check1_CheckInst_1_n15), .ZN(Check1_CheckInst_1_n96) );
  NOR2_X1 Check1_CheckInst_1_U14 ( .A1(Check1_CheckInst_1_n14), .A2(
        Check1_CheckInst_1_n13), .ZN(Check1_CheckInst_1_n15) );
  NAND2_X1 Check1_CheckInst_1_U13 ( .A1(Check1_CheckInst_1_n12), .A2(
        Check1_CheckInst_1_n11), .ZN(Check1_CheckInst_1_n13) );
  NOR2_X1 Check1_CheckInst_1_U12 ( .A1(Check1_CheckInst_1_n10), .A2(
        Check1_CheckInst_1_n9), .ZN(Check1_CheckInst_1_n11) );
  XOR2_X1 Check1_CheckInst_1_U11 ( .A(Red_MC_output[25]), .B(
        Red_SignaltoCheck[73]), .Z(Check1_CheckInst_1_n9) );
  XOR2_X1 Check1_CheckInst_1_U10 ( .A(Red_MC_output[37]), .B(
        Red_SignaltoCheck[85]), .Z(Check1_CheckInst_1_n10) );
  NOR2_X1 Check1_CheckInst_1_U9 ( .A1(Check1_CheckInst_1_n8), .A2(
        Check1_CheckInst_1_n7), .ZN(Check1_CheckInst_1_n12) );
  XOR2_X1 Check1_CheckInst_1_U8 ( .A(Red_MC_output[28]), .B(
        Red_SignaltoCheck[76]), .Z(Check1_CheckInst_1_n7) );
  XOR2_X1 Check1_CheckInst_1_U7 ( .A(Red_MC_output[22]), .B(
        Red_SignaltoCheck[70]), .Z(Check1_CheckInst_1_n8) );
  NAND2_X1 Check1_CheckInst_1_U6 ( .A1(Check1_CheckInst_1_n6), .A2(
        Check1_CheckInst_1_n5), .ZN(Check1_CheckInst_1_n14) );
  XNOR2_X1 Check1_CheckInst_1_U5 ( .A(Red_ShiftRowsOutput[37]), .B(
        Red_SignaltoCheck[133]), .ZN(Check1_CheckInst_1_n5) );
  XNOR2_X1 Check1_CheckInst_1_U4 ( .A(Red_ShiftRowsOutput[40]), .B(
        Red_SignaltoCheck[136]), .ZN(Check1_CheckInst_1_n6) );
  NOR2_X1 Check1_CheckInst_1_U3 ( .A1(Check1_CheckInst_1_n4), .A2(
        Check1_CheckInst_1_n3), .ZN(Check1_CheckInst_1_n16) );
  XOR2_X1 Check1_CheckInst_1_U2 ( .A(Red_ShiftRowsOutput[31]), .B(
        Red_SignaltoCheck[127]), .Z(Check1_CheckInst_1_n3) );
  XOR2_X1 Check1_CheckInst_1_U1 ( .A(Red_ShiftRowsOutput[43]), .B(
        Red_SignaltoCheck[139]), .Z(Check1_CheckInst_1_n4) );
  NOR2_X1 Check1_CheckInst_2_U95 ( .A1(Check1_CheckInst_2_n96), .A2(
        Check1_CheckInst_2_n95), .ZN(Error[2]) );
  NAND2_X1 Check1_CheckInst_2_U94 ( .A1(Check1_CheckInst_2_n94), .A2(
        Check1_CheckInst_2_n93), .ZN(Check1_CheckInst_2_n95) );
  NOR2_X1 Check1_CheckInst_2_U93 ( .A1(Check1_CheckInst_2_n92), .A2(
        Check1_CheckInst_2_n91), .ZN(Check1_CheckInst_2_n93) );
  NAND2_X1 Check1_CheckInst_2_U92 ( .A1(Check1_CheckInst_2_n90), .A2(
        Check1_CheckInst_2_n89), .ZN(Check1_CheckInst_2_n91) );
  NOR2_X1 Check1_CheckInst_2_U91 ( .A1(Check1_CheckInst_2_n88), .A2(
        Check1_CheckInst_2_n87), .ZN(Check1_CheckInst_2_n89) );
  NAND2_X1 Check1_CheckInst_2_U90 ( .A1(Check1_CheckInst_2_n86), .A2(
        Check1_CheckInst_2_n85), .ZN(Check1_CheckInst_2_n87) );
  NOR2_X1 Check1_CheckInst_2_U89 ( .A1(Check1_CheckInst_2_n84), .A2(
        Check1_CheckInst_2_n83), .ZN(Check1_CheckInst_2_n85) );
  XOR2_X1 Check1_CheckInst_2_U88 ( .A(Red_AddRoundKeyOutput[23]), .B(
        Red_SignaltoCheck[23]), .Z(Check1_CheckInst_2_n83) );
  XOR2_X1 Check1_CheckInst_2_U87 ( .A(Red_AddRoundKeyOutput[17]), .B(
        Red_SignaltoCheck[17]), .Z(Check1_CheckInst_2_n84) );
  XNOR2_X1 Check1_CheckInst_2_U86 ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[11]), .ZN(Check1_CheckInst_2_n86) );
  NAND2_X1 Check1_CheckInst_2_U85 ( .A1(Check1_CheckInst_2_n82), .A2(
        Check1_CheckInst_2_n81), .ZN(Check1_CheckInst_2_n88) );
  NOR2_X1 Check1_CheckInst_2_U84 ( .A1(Check1_CheckInst_2_n80), .A2(
        Check1_CheckInst_2_n79), .ZN(Check1_CheckInst_2_n81) );
  NAND2_X1 Check1_CheckInst_2_U83 ( .A1(Check1_CheckInst_2_n78), .A2(
        Check1_CheckInst_2_n77), .ZN(Check1_CheckInst_2_n79) );
  NOR2_X1 Check1_CheckInst_2_U82 ( .A1(Check1_CheckInst_2_n76), .A2(
        Check1_CheckInst_2_n75), .ZN(Check1_CheckInst_2_n77) );
  XOR2_X1 Check1_CheckInst_2_U81 ( .A(Red_AddRoundKeyOutput[26]), .B(
        Red_SignaltoCheck[26]), .Z(Check1_CheckInst_2_n75) );
  XOR2_X1 Check1_CheckInst_2_U80 ( .A(Red_AddRoundKeyOutput[29]), .B(
        Red_SignaltoCheck[29]), .Z(Check1_CheckInst_2_n76) );
  XNOR2_X1 Check1_CheckInst_2_U79 ( .A(Red_AddRoundKeyOutput[32]), .B(
        Red_SignaltoCheck[32]), .ZN(Check1_CheckInst_2_n78) );
  NAND2_X1 Check1_CheckInst_2_U78 ( .A1(Check1_CheckInst_2_n74), .A2(
        Check1_CheckInst_2_n73), .ZN(Check1_CheckInst_2_n80) );
  NOR2_X1 Check1_CheckInst_2_U77 ( .A1(Check1_CheckInst_2_n72), .A2(
        Check1_CheckInst_2_n71), .ZN(Check1_CheckInst_2_n73) );
  NAND2_X1 Check1_CheckInst_2_U76 ( .A1(Check1_CheckInst_2_n70), .A2(
        Check1_CheckInst_2_n69), .ZN(Check1_CheckInst_2_n71) );
  NOR2_X1 Check1_CheckInst_2_U75 ( .A1(Check1_CheckInst_2_n68), .A2(
        Check1_CheckInst_2_n67), .ZN(Check1_CheckInst_2_n69) );
  XOR2_X1 Check1_CheckInst_2_U74 ( .A(Red_ShiftRowsOutput[26]), .B(
        Red_SignaltoCheck[122]), .Z(Check1_CheckInst_2_n68) );
  XNOR2_X1 Check1_CheckInst_2_U73 ( .A(Red_ShiftRowsOutput[11]), .B(
        Red_SignaltoCheck[107]), .ZN(Check1_CheckInst_2_n70) );
  NAND2_X1 Check1_CheckInst_2_U72 ( .A1(Check1_CheckInst_2_n66), .A2(
        Check1_CheckInst_2_n65), .ZN(Check1_CheckInst_2_n72) );
  NOR2_X1 Check1_CheckInst_2_U71 ( .A1(Check1_CheckInst_2_n64), .A2(
        Check1_CheckInst_2_n63), .ZN(Check1_CheckInst_2_n65) );
  NOR2_X1 Check1_CheckInst_2_U70 ( .A1(Check1_CheckInst_2_n62), .A2(
        Check1_CheckInst_2_n61), .ZN(Check1_CheckInst_2_n66) );
  XNOR2_X1 Check1_CheckInst_2_U69 ( .A(Red_SignaltoCheck[113]), .B(
        Red_ShiftRowsOutput[17]), .ZN(Check1_CheckInst_2_n74) );
  XNOR2_X1 Check1_CheckInst_2_U68 ( .A(Red_SignaltoCheck[20]), .B(
        Red_AddRoundKeyOutput[20]), .ZN(Check1_CheckInst_2_n82) );
  XNOR2_X1 Check1_CheckInst_2_U67 ( .A(Red_SignaltoCheck[8]), .B(
        Red_AddRoundKeyOutput[8]), .ZN(Check1_CheckInst_2_n90) );
  NAND2_X1 Check1_CheckInst_2_U66 ( .A1(Check1_CheckInst_2_n60), .A2(
        Check1_CheckInst_2_n59), .ZN(Check1_CheckInst_2_n92) );
  NOR2_X1 Check1_CheckInst_2_U65 ( .A1(Check1_CheckInst_2_n58), .A2(
        Check1_CheckInst_2_n57), .ZN(Check1_CheckInst_2_n59) );
  NAND2_X1 Check1_CheckInst_2_U64 ( .A1(Check1_CheckInst_2_n56), .A2(
        Check1_CheckInst_2_n55), .ZN(Check1_CheckInst_2_n57) );
  NOR2_X1 Check1_CheckInst_2_U63 ( .A1(Check1_CheckInst_2_n54), .A2(
        Check1_CheckInst_2_n53), .ZN(Check1_CheckInst_2_n55) );
  XOR2_X1 Check1_CheckInst_2_U62 ( .A(Red_AddRoundKeyOutput[38]), .B(
        Red_SignaltoCheck[38]), .Z(Check1_CheckInst_2_n53) );
  XOR2_X1 Check1_CheckInst_2_U61 ( .A(Red_MC_output[2]), .B(
        Red_SignaltoCheck[50]), .Z(Check1_CheckInst_2_n54) );
  XNOR2_X1 Check1_CheckInst_2_U60 ( .A(Red_AddRoundKeyOutput[35]), .B(
        Red_SignaltoCheck[35]), .ZN(Check1_CheckInst_2_n56) );
  NAND2_X1 Check1_CheckInst_2_U59 ( .A1(Check1_CheckInst_2_n52), .A2(
        Check1_CheckInst_2_n51), .ZN(Check1_CheckInst_2_n58) );
  NOR2_X1 Check1_CheckInst_2_U58 ( .A1(Check1_CheckInst_2_n50), .A2(
        Check1_CheckInst_2_n49), .ZN(Check1_CheckInst_2_n51) );
  NAND2_X1 Check1_CheckInst_2_U57 ( .A1(Check1_CheckInst_2_n48), .A2(
        Check1_CheckInst_2_n47), .ZN(Check1_CheckInst_2_n49) );
  NOR2_X1 Check1_CheckInst_2_U56 ( .A1(Check1_CheckInst_2_n46), .A2(
        Check1_CheckInst_2_n45), .ZN(Check1_CheckInst_2_n47) );
  XOR2_X1 Check1_CheckInst_2_U55 ( .A(Red_MC_output[11]), .B(
        Red_SignaltoCheck[59]), .Z(Check1_CheckInst_2_n45) );
  XOR2_X1 Check1_CheckInst_2_U54 ( .A(Red_MC_output[5]), .B(
        Red_SignaltoCheck[53]), .Z(Check1_CheckInst_2_n46) );
  XNOR2_X1 Check1_CheckInst_2_U53 ( .A(Red_AddRoundKeyOutput[47]), .B(
        Red_SignaltoCheck[47]), .ZN(Check1_CheckInst_2_n48) );
  NAND2_X1 Check1_CheckInst_2_U52 ( .A1(Check1_CheckInst_2_n44), .A2(
        Check1_CheckInst_2_n43), .ZN(Check1_CheckInst_2_n50) );
  NOR2_X1 Check1_CheckInst_2_U51 ( .A1(Check1_CheckInst_2_n42), .A2(
        Check1_CheckInst_2_n41), .ZN(Check1_CheckInst_2_n43) );
  NAND2_X1 Check1_CheckInst_2_U50 ( .A1(Check1_CheckInst_2_n40), .A2(
        Check1_CheckInst_2_n39), .ZN(Check1_CheckInst_2_n41) );
  NOR2_X1 Check1_CheckInst_2_U49 ( .A1(Check1_CheckInst_2_n38), .A2(
        Check1_CheckInst_2_n37), .ZN(Check1_CheckInst_2_n39) );
  XOR2_X1 Check1_CheckInst_2_U48 ( .A(Red_MC_output[14]), .B(
        Red_SignaltoCheck[62]), .Z(Check1_CheckInst_2_n37) );
  XOR2_X1 Check1_CheckInst_2_U47 ( .A(Red_MC_output[17]), .B(
        Red_SignaltoCheck[65]), .Z(Check1_CheckInst_2_n38) );
  XNOR2_X1 Check1_CheckInst_2_U46 ( .A(Red_MC_output[20]), .B(
        Red_SignaltoCheck[68]), .ZN(Check1_CheckInst_2_n40) );
  NAND2_X1 Check1_CheckInst_2_U45 ( .A1(Check1_CheckInst_2_n36), .A2(
        Check1_CheckInst_2_n35), .ZN(Check1_CheckInst_2_n42) );
  NOR2_X1 Check1_CheckInst_2_U44 ( .A1(Check1_CheckInst_2_n34), .A2(
        Check1_CheckInst_2_n33), .ZN(Check1_CheckInst_2_n35) );
  XOR2_X1 Check1_CheckInst_2_U43 ( .A(Red_ShiftRowsOutput[47]), .B(
        Red_SignaltoCheck[143]), .Z(Check1_CheckInst_2_n33) );
  XOR2_X1 Check1_CheckInst_2_U42 ( .A(Red_SignaltoCheck[5]), .B(
        Red_AddRoundKeyOutput[5]), .Z(Check1_CheckInst_2_n34) );
  NOR2_X1 Check1_CheckInst_2_U41 ( .A1(Check1_CheckInst_2_n32), .A2(
        Check1_CheckInst_2_n31), .ZN(Check1_CheckInst_2_n36) );
  XOR2_X1 Check1_CheckInst_2_U40 ( .A(Red_AddRoundKeyOutput[2]), .B(
        Red_SignaltoCheck[2]), .Z(Check1_CheckInst_2_n31) );
  XOR2_X1 Check1_CheckInst_2_U39 ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[14]), .Z(Check1_CheckInst_2_n32) );
  XNOR2_X1 Check1_CheckInst_2_U38 ( .A(Red_SignaltoCheck[56]), .B(
        Red_MC_output[8]), .ZN(Check1_CheckInst_2_n44) );
  XNOR2_X1 Check1_CheckInst_2_U37 ( .A(Red_SignaltoCheck[44]), .B(
        Red_AddRoundKeyOutput[44]), .ZN(Check1_CheckInst_2_n52) );
  XNOR2_X1 Check1_CheckInst_2_U36 ( .A(Red_SignaltoCheck[41]), .B(
        Red_AddRoundKeyOutput[41]), .ZN(Check1_CheckInst_2_n60) );
  NOR2_X1 Check1_CheckInst_2_U35 ( .A1(Check1_CheckInst_2_n30), .A2(
        Check1_CheckInst_2_n29), .ZN(Check1_CheckInst_2_n94) );
  NAND2_X1 Check1_CheckInst_2_U34 ( .A1(Check1_CheckInst_2_n28), .A2(
        Check1_CheckInst_2_n27), .ZN(Check1_CheckInst_2_n29) );
  NOR2_X1 Check1_CheckInst_2_U33 ( .A1(Check1_CheckInst_2_n26), .A2(
        Check1_CheckInst_2_n25), .ZN(Check1_CheckInst_2_n27) );
  NAND2_X1 Check1_CheckInst_2_U32 ( .A1(Check1_CheckInst_2_n24), .A2(
        Check1_CheckInst_2_n23), .ZN(Check1_CheckInst_2_n25) );
  NAND2_X1 Check1_CheckInst_2_U31 ( .A1(Check1_CheckInst_2_n22), .A2(
        Check1_CheckInst_2_n21), .ZN(Check1_CheckInst_2_n26) );
  XNOR2_X1 Check1_CheckInst_2_U30 ( .A(Red_MC_output[44]), .B(
        Red_SignaltoCheck[92]), .ZN(Check1_CheckInst_2_n21) );
  NOR2_X1 Check1_CheckInst_2_U29 ( .A1(Check1_CheckInst_2_n20), .A2(
        Check1_CheckInst_2_n19), .ZN(Check1_CheckInst_2_n28) );
  XOR2_X1 Check1_CheckInst_2_U28 ( .A(Red_MC_output[47]), .B(
        Red_SignaltoCheck[95]), .Z(Check1_CheckInst_2_n19) );
  XOR2_X1 Check1_CheckInst_2_U27 ( .A(Red_MC_output[41]), .B(
        Red_SignaltoCheck[89]), .Z(Check1_CheckInst_2_n20) );
  NAND2_X1 Check1_CheckInst_2_U26 ( .A1(Check1_CheckInst_2_n18), .A2(
        Check1_CheckInst_2_n17), .ZN(Check1_CheckInst_2_n30) );
  XNOR2_X1 Check1_CheckInst_2_U25 ( .A(Red_MC_output[32]), .B(
        Red_SignaltoCheck[80]), .ZN(Check1_CheckInst_2_n17) );
  XNOR2_X1 Check1_CheckInst_2_U24 ( .A(Red_MC_output[35]), .B(
        Red_SignaltoCheck[83]), .ZN(Check1_CheckInst_2_n18) );
  NAND2_X1 Check1_CheckInst_2_U23 ( .A1(Check1_CheckInst_2_n16), .A2(
        Check1_CheckInst_2_n15), .ZN(Check1_CheckInst_2_n96) );
  NOR2_X1 Check1_CheckInst_2_U22 ( .A1(Check1_CheckInst_2_n14), .A2(
        Check1_CheckInst_2_n13), .ZN(Check1_CheckInst_2_n15) );
  NAND2_X1 Check1_CheckInst_2_U21 ( .A1(Check1_CheckInst_2_n12), .A2(
        Check1_CheckInst_2_n11), .ZN(Check1_CheckInst_2_n13) );
  NOR2_X1 Check1_CheckInst_2_U20 ( .A1(Check1_CheckInst_2_n10), .A2(
        Check1_CheckInst_2_n9), .ZN(Check1_CheckInst_2_n11) );
  XOR2_X1 Check1_CheckInst_2_U19 ( .A(Red_MC_output[26]), .B(
        Red_SignaltoCheck[74]), .Z(Check1_CheckInst_2_n9) );
  XOR2_X1 Check1_CheckInst_2_U18 ( .A(Red_MC_output[38]), .B(
        Red_SignaltoCheck[86]), .Z(Check1_CheckInst_2_n10) );
  NOR2_X1 Check1_CheckInst_2_U17 ( .A1(Check1_CheckInst_2_n8), .A2(
        Check1_CheckInst_2_n7), .ZN(Check1_CheckInst_2_n12) );
  XOR2_X1 Check1_CheckInst_2_U16 ( .A(Red_MC_output[29]), .B(
        Red_SignaltoCheck[77]), .Z(Check1_CheckInst_2_n7) );
  XOR2_X1 Check1_CheckInst_2_U15 ( .A(Red_MC_output[23]), .B(
        Red_SignaltoCheck[71]), .Z(Check1_CheckInst_2_n8) );
  NAND2_X1 Check1_CheckInst_2_U14 ( .A1(Check1_CheckInst_2_n6), .A2(
        Check1_CheckInst_2_n5), .ZN(Check1_CheckInst_2_n14) );
  XNOR2_X1 Check1_CheckInst_2_U13 ( .A(Red_ShiftRowsOutput[38]), .B(
        Red_SignaltoCheck[134]), .ZN(Check1_CheckInst_2_n5) );
  XNOR2_X1 Check1_CheckInst_2_U12 ( .A(Red_ShiftRowsOutput[41]), .B(
        Red_SignaltoCheck[137]), .ZN(Check1_CheckInst_2_n6) );
  NOR2_X1 Check1_CheckInst_2_U11 ( .A1(Check1_CheckInst_2_n4), .A2(
        Check1_CheckInst_2_n3), .ZN(Check1_CheckInst_2_n16) );
  XOR2_X1 Check1_CheckInst_2_U10 ( .A(Red_ShiftRowsOutput[44]), .B(
        Red_SignaltoCheck[140]), .Z(Check1_CheckInst_2_n4) );
  XOR2_X1 Check1_CheckInst_2_U9 ( .A(Red_ShiftRowsOutput[29]), .B(
        Red_SignaltoCheck[125]), .Z(Check1_CheckInst_2_n62) );
  XOR2_X1 Check1_CheckInst_2_U8 ( .A(Red_ShiftRowsOutput[32]), .B(
        Red_SignaltoCheck[128]), .Z(Check1_CheckInst_2_n3) );
  XOR2_X1 Check1_CheckInst_2_U7 ( .A(Red_ShiftRowsOutput[35]), .B(
        Red_SignaltoCheck[131]), .Z(Check1_CheckInst_2_n61) );
  XNOR2_X1 Check1_CheckInst_2_U6 ( .A(Red_ShiftRowsOutput[8]), .B(
        Red_SignaltoCheck[104]), .ZN(Check1_CheckInst_2_n22) );
  XOR2_X1 Check1_CheckInst_2_U5 ( .A(Red_ShiftRowsOutput[23]), .B(
        Red_SignaltoCheck[119]), .Z(Check1_CheckInst_2_n64) );
  XNOR2_X1 Check1_CheckInst_2_U4 ( .A(Red_ShiftRowsOutput[5]), .B(
        Red_SignaltoCheck[101]), .ZN(Check1_CheckInst_2_n24) );
  XOR2_X1 Check1_CheckInst_2_U3 ( .A(Red_ShiftRowsOutput[20]), .B(
        Red_SignaltoCheck[116]), .Z(Check1_CheckInst_2_n63) );
  XNOR2_X1 Check1_CheckInst_2_U2 ( .A(Red_ShiftRowsOutput[2]), .B(
        Red_SignaltoCheck[98]), .ZN(Check1_CheckInst_2_n23) );
  XOR2_X1 Check1_CheckInst_2_U1 ( .A(Red_ShiftRowsOutput[14]), .B(
        Red_SignaltoCheck[110]), .Z(Check1_CheckInst_2_n67) );
endmodule

