
module LED64Enc ( clk, Plaintext, Key, Ciphertext, ErrorFlag );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* fiver="clock" *)input clk;
  output ErrorFlag;
  wire   n4, SubCellInst_LFInst_0_LFInst_0_n9,
         SubCellInst_LFInst_0_LFInst_0_n8, SubCellInst_LFInst_0_LFInst_0_n7,
         SubCellInst_LFInst_0_LFInst_0_n10, SubCellInst_LFInst_0_LFInst_1_n26,
         SubCellInst_LFInst_0_LFInst_1_n25, SubCellInst_LFInst_0_LFInst_1_n24,
         SubCellInst_LFInst_0_LFInst_1_n23, SubCellInst_LFInst_0_LFInst_1_n22,
         SubCellInst_LFInst_0_LFInst_1_n21, SubCellInst_LFInst_0_LFInst_1_n20,
         SubCellInst_LFInst_0_LFInst_1_n19, SubCellInst_LFInst_0_LFInst_1_n18,
         SubCellInst_LFInst_0_LFInst_2_n28, SubCellInst_LFInst_0_LFInst_2_n27,
         SubCellInst_LFInst_0_LFInst_2_n26, SubCellInst_LFInst_0_LFInst_2_n25,
         SubCellInst_LFInst_0_LFInst_2_n24, SubCellInst_LFInst_0_LFInst_2_n23,
         SubCellInst_LFInst_0_LFInst_2_n22, SubCellInst_LFInst_0_LFInst_3_n26,
         SubCellInst_LFInst_0_LFInst_3_n25, SubCellInst_LFInst_0_LFInst_3_n24,
         SubCellInst_LFInst_0_LFInst_3_n23, SubCellInst_LFInst_0_LFInst_3_n22,
         SubCellInst_LFInst_0_LFInst_3_n21, SubCellInst_LFInst_0_LFInst_3_n20,
         SubCellInst_LFInst_0_LFInst_3_n19, SubCellInst_LFInst_1_LFInst_0_n9,
         SubCellInst_LFInst_1_LFInst_0_n8, SubCellInst_LFInst_1_LFInst_0_n7,
         SubCellInst_LFInst_1_LFInst_0_n10, SubCellInst_LFInst_1_LFInst_1_n26,
         SubCellInst_LFInst_1_LFInst_1_n25, SubCellInst_LFInst_1_LFInst_1_n24,
         SubCellInst_LFInst_1_LFInst_1_n23, SubCellInst_LFInst_1_LFInst_1_n22,
         SubCellInst_LFInst_1_LFInst_1_n21, SubCellInst_LFInst_1_LFInst_1_n20,
         SubCellInst_LFInst_1_LFInst_1_n19, SubCellInst_LFInst_1_LFInst_1_n18,
         SubCellInst_LFInst_1_LFInst_2_n28, SubCellInst_LFInst_1_LFInst_2_n27,
         SubCellInst_LFInst_1_LFInst_2_n26, SubCellInst_LFInst_1_LFInst_2_n25,
         SubCellInst_LFInst_1_LFInst_2_n24, SubCellInst_LFInst_1_LFInst_2_n23,
         SubCellInst_LFInst_1_LFInst_2_n22, SubCellInst_LFInst_1_LFInst_3_n26,
         SubCellInst_LFInst_1_LFInst_3_n25, SubCellInst_LFInst_1_LFInst_3_n24,
         SubCellInst_LFInst_1_LFInst_3_n23, SubCellInst_LFInst_1_LFInst_3_n22,
         SubCellInst_LFInst_1_LFInst_3_n21, SubCellInst_LFInst_1_LFInst_3_n20,
         SubCellInst_LFInst_1_LFInst_3_n19, SubCellInst_LFInst_2_LFInst_0_n9,
         SubCellInst_LFInst_2_LFInst_0_n8, SubCellInst_LFInst_2_LFInst_0_n7,
         SubCellInst_LFInst_2_LFInst_0_n10, SubCellInst_LFInst_2_LFInst_1_n26,
         SubCellInst_LFInst_2_LFInst_1_n25, SubCellInst_LFInst_2_LFInst_1_n24,
         SubCellInst_LFInst_2_LFInst_1_n23, SubCellInst_LFInst_2_LFInst_1_n22,
         SubCellInst_LFInst_2_LFInst_1_n21, SubCellInst_LFInst_2_LFInst_1_n20,
         SubCellInst_LFInst_2_LFInst_1_n19, SubCellInst_LFInst_2_LFInst_1_n18,
         SubCellInst_LFInst_2_LFInst_2_n28, SubCellInst_LFInst_2_LFInst_2_n27,
         SubCellInst_LFInst_2_LFInst_2_n26, SubCellInst_LFInst_2_LFInst_2_n25,
         SubCellInst_LFInst_2_LFInst_2_n24, SubCellInst_LFInst_2_LFInst_2_n23,
         SubCellInst_LFInst_2_LFInst_2_n22, SubCellInst_LFInst_2_LFInst_3_n26,
         SubCellInst_LFInst_2_LFInst_3_n25, SubCellInst_LFInst_2_LFInst_3_n24,
         SubCellInst_LFInst_2_LFInst_3_n23, SubCellInst_LFInst_2_LFInst_3_n22,
         SubCellInst_LFInst_2_LFInst_3_n21, SubCellInst_LFInst_2_LFInst_3_n20,
         SubCellInst_LFInst_2_LFInst_3_n19, SubCellInst_LFInst_3_LFInst_0_n9,
         SubCellInst_LFInst_3_LFInst_0_n8, SubCellInst_LFInst_3_LFInst_0_n7,
         SubCellInst_LFInst_3_LFInst_0_n10, SubCellInst_LFInst_3_LFInst_1_n26,
         SubCellInst_LFInst_3_LFInst_1_n25, SubCellInst_LFInst_3_LFInst_1_n24,
         SubCellInst_LFInst_3_LFInst_1_n23, SubCellInst_LFInst_3_LFInst_1_n22,
         SubCellInst_LFInst_3_LFInst_1_n21, SubCellInst_LFInst_3_LFInst_1_n20,
         SubCellInst_LFInst_3_LFInst_1_n19, SubCellInst_LFInst_3_LFInst_1_n18,
         SubCellInst_LFInst_3_LFInst_2_n28, SubCellInst_LFInst_3_LFInst_2_n27,
         SubCellInst_LFInst_3_LFInst_2_n26, SubCellInst_LFInst_3_LFInst_2_n25,
         SubCellInst_LFInst_3_LFInst_2_n24, SubCellInst_LFInst_3_LFInst_2_n23,
         SubCellInst_LFInst_3_LFInst_2_n22, SubCellInst_LFInst_3_LFInst_3_n26,
         SubCellInst_LFInst_3_LFInst_3_n25, SubCellInst_LFInst_3_LFInst_3_n24,
         SubCellInst_LFInst_3_LFInst_3_n23, SubCellInst_LFInst_3_LFInst_3_n22,
         SubCellInst_LFInst_3_LFInst_3_n21, SubCellInst_LFInst_3_LFInst_3_n20,
         SubCellInst_LFInst_3_LFInst_3_n19, SubCellInst_LFInst_4_LFInst_0_n8,
         SubCellInst_LFInst_4_LFInst_0_n7, SubCellInst_LFInst_4_LFInst_0_n6,
         SubCellInst_LFInst_4_LFInst_1_n26, SubCellInst_LFInst_4_LFInst_1_n25,
         SubCellInst_LFInst_4_LFInst_1_n24, SubCellInst_LFInst_4_LFInst_1_n23,
         SubCellInst_LFInst_4_LFInst_1_n22, SubCellInst_LFInst_4_LFInst_1_n21,
         SubCellInst_LFInst_4_LFInst_1_n20, SubCellInst_LFInst_4_LFInst_1_n19,
         SubCellInst_LFInst_4_LFInst_1_n18, SubCellInst_LFInst_4_LFInst_2_n29,
         SubCellInst_LFInst_4_LFInst_2_n28, SubCellInst_LFInst_4_LFInst_2_n27,
         SubCellInst_LFInst_4_LFInst_2_n26, SubCellInst_LFInst_4_LFInst_2_n25,
         SubCellInst_LFInst_4_LFInst_2_n24, SubCellInst_LFInst_4_LFInst_2_n23,
         SubCellInst_LFInst_4_LFInst_2_n22, SubCellInst_LFInst_4_LFInst_3_n26,
         SubCellInst_LFInst_4_LFInst_3_n25, SubCellInst_LFInst_4_LFInst_3_n24,
         SubCellInst_LFInst_4_LFInst_3_n23, SubCellInst_LFInst_4_LFInst_3_n22,
         SubCellInst_LFInst_4_LFInst_3_n21, SubCellInst_LFInst_4_LFInst_3_n20,
         SubCellInst_LFInst_4_LFInst_3_n19, SubCellInst_LFInst_5_LFInst_0_n8,
         SubCellInst_LFInst_5_LFInst_0_n7, SubCellInst_LFInst_5_LFInst_0_n6,
         SubCellInst_LFInst_5_LFInst_1_n26, SubCellInst_LFInst_5_LFInst_1_n25,
         SubCellInst_LFInst_5_LFInst_1_n24, SubCellInst_LFInst_5_LFInst_1_n23,
         SubCellInst_LFInst_5_LFInst_1_n22, SubCellInst_LFInst_5_LFInst_1_n21,
         SubCellInst_LFInst_5_LFInst_1_n20, SubCellInst_LFInst_5_LFInst_1_n19,
         SubCellInst_LFInst_5_LFInst_1_n18, SubCellInst_LFInst_5_LFInst_2_n29,
         SubCellInst_LFInst_5_LFInst_2_n28, SubCellInst_LFInst_5_LFInst_2_n27,
         SubCellInst_LFInst_5_LFInst_2_n26, SubCellInst_LFInst_5_LFInst_2_n25,
         SubCellInst_LFInst_5_LFInst_2_n24, SubCellInst_LFInst_5_LFInst_2_n23,
         SubCellInst_LFInst_5_LFInst_2_n22, SubCellInst_LFInst_5_LFInst_3_n26,
         SubCellInst_LFInst_5_LFInst_3_n25, SubCellInst_LFInst_5_LFInst_3_n24,
         SubCellInst_LFInst_5_LFInst_3_n23, SubCellInst_LFInst_5_LFInst_3_n22,
         SubCellInst_LFInst_5_LFInst_3_n21, SubCellInst_LFInst_5_LFInst_3_n20,
         SubCellInst_LFInst_5_LFInst_3_n19, SubCellInst_LFInst_6_LFInst_0_n8,
         SubCellInst_LFInst_6_LFInst_0_n7, SubCellInst_LFInst_6_LFInst_0_n6,
         SubCellInst_LFInst_6_LFInst_1_n26, SubCellInst_LFInst_6_LFInst_1_n25,
         SubCellInst_LFInst_6_LFInst_1_n24, SubCellInst_LFInst_6_LFInst_1_n23,
         SubCellInst_LFInst_6_LFInst_1_n22, SubCellInst_LFInst_6_LFInst_1_n21,
         SubCellInst_LFInst_6_LFInst_1_n20, SubCellInst_LFInst_6_LFInst_1_n19,
         SubCellInst_LFInst_6_LFInst_1_n18, SubCellInst_LFInst_6_LFInst_2_n29,
         SubCellInst_LFInst_6_LFInst_2_n28, SubCellInst_LFInst_6_LFInst_2_n27,
         SubCellInst_LFInst_6_LFInst_2_n26, SubCellInst_LFInst_6_LFInst_2_n25,
         SubCellInst_LFInst_6_LFInst_2_n24, SubCellInst_LFInst_6_LFInst_2_n23,
         SubCellInst_LFInst_6_LFInst_2_n22, SubCellInst_LFInst_6_LFInst_3_n26,
         SubCellInst_LFInst_6_LFInst_3_n25, SubCellInst_LFInst_6_LFInst_3_n24,
         SubCellInst_LFInst_6_LFInst_3_n23, SubCellInst_LFInst_6_LFInst_3_n22,
         SubCellInst_LFInst_6_LFInst_3_n21, SubCellInst_LFInst_6_LFInst_3_n20,
         SubCellInst_LFInst_6_LFInst_3_n19, SubCellInst_LFInst_7_LFInst_0_n8,
         SubCellInst_LFInst_7_LFInst_0_n7, SubCellInst_LFInst_7_LFInst_0_n6,
         SubCellInst_LFInst_7_LFInst_1_n26, SubCellInst_LFInst_7_LFInst_1_n25,
         SubCellInst_LFInst_7_LFInst_1_n24, SubCellInst_LFInst_7_LFInst_1_n23,
         SubCellInst_LFInst_7_LFInst_1_n22, SubCellInst_LFInst_7_LFInst_1_n21,
         SubCellInst_LFInst_7_LFInst_1_n20, SubCellInst_LFInst_7_LFInst_1_n19,
         SubCellInst_LFInst_7_LFInst_1_n18, SubCellInst_LFInst_7_LFInst_2_n29,
         SubCellInst_LFInst_7_LFInst_2_n28, SubCellInst_LFInst_7_LFInst_2_n27,
         SubCellInst_LFInst_7_LFInst_2_n26, SubCellInst_LFInst_7_LFInst_2_n25,
         SubCellInst_LFInst_7_LFInst_2_n24, SubCellInst_LFInst_7_LFInst_2_n23,
         SubCellInst_LFInst_7_LFInst_2_n22, SubCellInst_LFInst_7_LFInst_3_n26,
         SubCellInst_LFInst_7_LFInst_3_n25, SubCellInst_LFInst_7_LFInst_3_n24,
         SubCellInst_LFInst_7_LFInst_3_n23, SubCellInst_LFInst_7_LFInst_3_n22,
         SubCellInst_LFInst_7_LFInst_3_n21, SubCellInst_LFInst_7_LFInst_3_n20,
         SubCellInst_LFInst_7_LFInst_3_n19, SubCellInst_LFInst_8_LFInst_0_n11,
         SubCellInst_LFInst_8_LFInst_0_n10, SubCellInst_LFInst_8_LFInst_0_n9,
         SubCellInst_LFInst_8_LFInst_0_n12, SubCellInst_LFInst_8_LFInst_1_n26,
         SubCellInst_LFInst_8_LFInst_1_n25, SubCellInst_LFInst_8_LFInst_1_n24,
         SubCellInst_LFInst_8_LFInst_1_n23, SubCellInst_LFInst_8_LFInst_1_n22,
         SubCellInst_LFInst_8_LFInst_1_n21, SubCellInst_LFInst_8_LFInst_1_n20,
         SubCellInst_LFInst_8_LFInst_1_n19, SubCellInst_LFInst_8_LFInst_1_n18,
         SubCellInst_LFInst_8_LFInst_2_n28, SubCellInst_LFInst_8_LFInst_2_n27,
         SubCellInst_LFInst_8_LFInst_2_n26, SubCellInst_LFInst_8_LFInst_2_n25,
         SubCellInst_LFInst_8_LFInst_2_n24, SubCellInst_LFInst_8_LFInst_2_n23,
         SubCellInst_LFInst_8_LFInst_2_n22, SubCellInst_LFInst_8_LFInst_3_n26,
         SubCellInst_LFInst_8_LFInst_3_n25, SubCellInst_LFInst_8_LFInst_3_n24,
         SubCellInst_LFInst_8_LFInst_3_n23, SubCellInst_LFInst_8_LFInst_3_n22,
         SubCellInst_LFInst_8_LFInst_3_n21, SubCellInst_LFInst_8_LFInst_3_n20,
         SubCellInst_LFInst_8_LFInst_3_n19, SubCellInst_LFInst_9_LFInst_0_n12,
         SubCellInst_LFInst_9_LFInst_0_n11, SubCellInst_LFInst_9_LFInst_0_n10,
         SubCellInst_LFInst_9_LFInst_0_n9, SubCellInst_LFInst_9_LFInst_1_n26,
         SubCellInst_LFInst_9_LFInst_1_n25, SubCellInst_LFInst_9_LFInst_1_n24,
         SubCellInst_LFInst_9_LFInst_1_n23, SubCellInst_LFInst_9_LFInst_1_n22,
         SubCellInst_LFInst_9_LFInst_1_n21, SubCellInst_LFInst_9_LFInst_1_n20,
         SubCellInst_LFInst_9_LFInst_1_n19, SubCellInst_LFInst_9_LFInst_1_n18,
         SubCellInst_LFInst_9_LFInst_2_n28, SubCellInst_LFInst_9_LFInst_2_n27,
         SubCellInst_LFInst_9_LFInst_2_n26, SubCellInst_LFInst_9_LFInst_2_n25,
         SubCellInst_LFInst_9_LFInst_2_n24, SubCellInst_LFInst_9_LFInst_2_n23,
         SubCellInst_LFInst_9_LFInst_2_n22, SubCellInst_LFInst_9_LFInst_3_n26,
         SubCellInst_LFInst_9_LFInst_3_n25, SubCellInst_LFInst_9_LFInst_3_n24,
         SubCellInst_LFInst_9_LFInst_3_n23, SubCellInst_LFInst_9_LFInst_3_n22,
         SubCellInst_LFInst_9_LFInst_3_n21, SubCellInst_LFInst_9_LFInst_3_n20,
         SubCellInst_LFInst_9_LFInst_3_n19, SubCellInst_LFInst_10_LFInst_0_n12,
         SubCellInst_LFInst_10_LFInst_0_n11,
         SubCellInst_LFInst_10_LFInst_0_n10, SubCellInst_LFInst_10_LFInst_0_n9,
         SubCellInst_LFInst_10_LFInst_1_n26,
         SubCellInst_LFInst_10_LFInst_1_n25,
         SubCellInst_LFInst_10_LFInst_1_n24,
         SubCellInst_LFInst_10_LFInst_1_n23,
         SubCellInst_LFInst_10_LFInst_1_n22,
         SubCellInst_LFInst_10_LFInst_1_n21,
         SubCellInst_LFInst_10_LFInst_1_n20,
         SubCellInst_LFInst_10_LFInst_1_n19,
         SubCellInst_LFInst_10_LFInst_1_n18,
         SubCellInst_LFInst_10_LFInst_2_n28,
         SubCellInst_LFInst_10_LFInst_2_n27,
         SubCellInst_LFInst_10_LFInst_2_n26,
         SubCellInst_LFInst_10_LFInst_2_n25,
         SubCellInst_LFInst_10_LFInst_2_n24,
         SubCellInst_LFInst_10_LFInst_2_n23,
         SubCellInst_LFInst_10_LFInst_2_n22,
         SubCellInst_LFInst_10_LFInst_3_n26,
         SubCellInst_LFInst_10_LFInst_3_n25,
         SubCellInst_LFInst_10_LFInst_3_n24,
         SubCellInst_LFInst_10_LFInst_3_n23,
         SubCellInst_LFInst_10_LFInst_3_n22,
         SubCellInst_LFInst_10_LFInst_3_n21,
         SubCellInst_LFInst_10_LFInst_3_n20,
         SubCellInst_LFInst_10_LFInst_3_n19,
         SubCellInst_LFInst_11_LFInst_0_n12,
         SubCellInst_LFInst_11_LFInst_0_n11,
         SubCellInst_LFInst_11_LFInst_0_n10, SubCellInst_LFInst_11_LFInst_0_n9,
         SubCellInst_LFInst_11_LFInst_1_n26,
         SubCellInst_LFInst_11_LFInst_1_n25,
         SubCellInst_LFInst_11_LFInst_1_n24,
         SubCellInst_LFInst_11_LFInst_1_n23,
         SubCellInst_LFInst_11_LFInst_1_n22,
         SubCellInst_LFInst_11_LFInst_1_n21,
         SubCellInst_LFInst_11_LFInst_1_n20,
         SubCellInst_LFInst_11_LFInst_1_n19,
         SubCellInst_LFInst_11_LFInst_1_n18,
         SubCellInst_LFInst_11_LFInst_2_n28,
         SubCellInst_LFInst_11_LFInst_2_n27,
         SubCellInst_LFInst_11_LFInst_2_n26,
         SubCellInst_LFInst_11_LFInst_2_n25,
         SubCellInst_LFInst_11_LFInst_2_n24,
         SubCellInst_LFInst_11_LFInst_2_n23,
         SubCellInst_LFInst_11_LFInst_2_n22,
         SubCellInst_LFInst_11_LFInst_3_n26,
         SubCellInst_LFInst_11_LFInst_3_n25,
         SubCellInst_LFInst_11_LFInst_3_n24,
         SubCellInst_LFInst_11_LFInst_3_n23,
         SubCellInst_LFInst_11_LFInst_3_n22,
         SubCellInst_LFInst_11_LFInst_3_n21,
         SubCellInst_LFInst_11_LFInst_3_n20,
         SubCellInst_LFInst_11_LFInst_3_n19, SubCellInst_LFInst_12_LFInst_0_n8,
         SubCellInst_LFInst_12_LFInst_0_n7, SubCellInst_LFInst_12_LFInst_0_n6,
         SubCellInst_LFInst_12_LFInst_0_n9, SubCellInst_LFInst_12_LFInst_1_n26,
         SubCellInst_LFInst_12_LFInst_1_n25,
         SubCellInst_LFInst_12_LFInst_1_n24,
         SubCellInst_LFInst_12_LFInst_1_n23,
         SubCellInst_LFInst_12_LFInst_1_n22,
         SubCellInst_LFInst_12_LFInst_1_n21,
         SubCellInst_LFInst_12_LFInst_1_n20,
         SubCellInst_LFInst_12_LFInst_1_n19,
         SubCellInst_LFInst_12_LFInst_1_n18,
         SubCellInst_LFInst_12_LFInst_2_n28,
         SubCellInst_LFInst_12_LFInst_2_n27,
         SubCellInst_LFInst_12_LFInst_2_n26,
         SubCellInst_LFInst_12_LFInst_2_n25,
         SubCellInst_LFInst_12_LFInst_2_n24,
         SubCellInst_LFInst_12_LFInst_2_n23,
         SubCellInst_LFInst_12_LFInst_2_n22,
         SubCellInst_LFInst_12_LFInst_3_n26,
         SubCellInst_LFInst_12_LFInst_3_n25,
         SubCellInst_LFInst_12_LFInst_3_n24,
         SubCellInst_LFInst_12_LFInst_3_n23,
         SubCellInst_LFInst_12_LFInst_3_n22,
         SubCellInst_LFInst_12_LFInst_3_n21,
         SubCellInst_LFInst_12_LFInst_3_n20,
         SubCellInst_LFInst_12_LFInst_3_n19, SubCellInst_LFInst_13_LFInst_0_n8,
         SubCellInst_LFInst_13_LFInst_0_n7, SubCellInst_LFInst_13_LFInst_0_n6,
         SubCellInst_LFInst_13_LFInst_0_n9, SubCellInst_LFInst_13_LFInst_1_n26,
         SubCellInst_LFInst_13_LFInst_1_n25,
         SubCellInst_LFInst_13_LFInst_1_n24,
         SubCellInst_LFInst_13_LFInst_1_n23,
         SubCellInst_LFInst_13_LFInst_1_n22,
         SubCellInst_LFInst_13_LFInst_1_n21,
         SubCellInst_LFInst_13_LFInst_1_n20,
         SubCellInst_LFInst_13_LFInst_1_n19,
         SubCellInst_LFInst_13_LFInst_1_n18,
         SubCellInst_LFInst_13_LFInst_2_n28,
         SubCellInst_LFInst_13_LFInst_2_n27,
         SubCellInst_LFInst_13_LFInst_2_n26,
         SubCellInst_LFInst_13_LFInst_2_n25,
         SubCellInst_LFInst_13_LFInst_2_n24,
         SubCellInst_LFInst_13_LFInst_2_n23,
         SubCellInst_LFInst_13_LFInst_2_n22,
         SubCellInst_LFInst_13_LFInst_3_n26,
         SubCellInst_LFInst_13_LFInst_3_n25,
         SubCellInst_LFInst_13_LFInst_3_n24,
         SubCellInst_LFInst_13_LFInst_3_n23,
         SubCellInst_LFInst_13_LFInst_3_n22,
         SubCellInst_LFInst_13_LFInst_3_n21,
         SubCellInst_LFInst_13_LFInst_3_n20,
         SubCellInst_LFInst_13_LFInst_3_n19, SubCellInst_LFInst_14_LFInst_0_n8,
         SubCellInst_LFInst_14_LFInst_0_n7, SubCellInst_LFInst_14_LFInst_0_n6,
         SubCellInst_LFInst_14_LFInst_0_n9, SubCellInst_LFInst_14_LFInst_1_n26,
         SubCellInst_LFInst_14_LFInst_1_n25,
         SubCellInst_LFInst_14_LFInst_1_n24,
         SubCellInst_LFInst_14_LFInst_1_n23,
         SubCellInst_LFInst_14_LFInst_1_n22,
         SubCellInst_LFInst_14_LFInst_1_n21,
         SubCellInst_LFInst_14_LFInst_1_n20,
         SubCellInst_LFInst_14_LFInst_1_n19,
         SubCellInst_LFInst_14_LFInst_1_n18,
         SubCellInst_LFInst_14_LFInst_2_n28,
         SubCellInst_LFInst_14_LFInst_2_n27,
         SubCellInst_LFInst_14_LFInst_2_n26,
         SubCellInst_LFInst_14_LFInst_2_n25,
         SubCellInst_LFInst_14_LFInst_2_n24,
         SubCellInst_LFInst_14_LFInst_2_n23,
         SubCellInst_LFInst_14_LFInst_2_n22,
         SubCellInst_LFInst_14_LFInst_3_n26,
         SubCellInst_LFInst_14_LFInst_3_n25,
         SubCellInst_LFInst_14_LFInst_3_n24,
         SubCellInst_LFInst_14_LFInst_3_n23,
         SubCellInst_LFInst_14_LFInst_3_n22,
         SubCellInst_LFInst_14_LFInst_3_n21,
         SubCellInst_LFInst_14_LFInst_3_n20,
         SubCellInst_LFInst_14_LFInst_3_n19, SubCellInst_LFInst_15_LFInst_0_n8,
         SubCellInst_LFInst_15_LFInst_0_n7, SubCellInst_LFInst_15_LFInst_0_n6,
         SubCellInst_LFInst_15_LFInst_0_n9, SubCellInst_LFInst_15_LFInst_1_n26,
         SubCellInst_LFInst_15_LFInst_1_n25,
         SubCellInst_LFInst_15_LFInst_1_n24,
         SubCellInst_LFInst_15_LFInst_1_n23,
         SubCellInst_LFInst_15_LFInst_1_n22,
         SubCellInst_LFInst_15_LFInst_1_n21,
         SubCellInst_LFInst_15_LFInst_1_n20,
         SubCellInst_LFInst_15_LFInst_1_n19,
         SubCellInst_LFInst_15_LFInst_1_n18,
         SubCellInst_LFInst_15_LFInst_2_n28,
         SubCellInst_LFInst_15_LFInst_2_n27,
         SubCellInst_LFInst_15_LFInst_2_n26,
         SubCellInst_LFInst_15_LFInst_2_n25,
         SubCellInst_LFInst_15_LFInst_2_n24,
         SubCellInst_LFInst_15_LFInst_2_n23,
         SubCellInst_LFInst_15_LFInst_2_n22,
         SubCellInst_LFInst_15_LFInst_3_n26,
         SubCellInst_LFInst_15_LFInst_3_n25,
         SubCellInst_LFInst_15_LFInst_3_n24,
         SubCellInst_LFInst_15_LFInst_3_n23,
         SubCellInst_LFInst_15_LFInst_3_n22,
         SubCellInst_LFInst_15_LFInst_3_n21,
         SubCellInst_LFInst_15_LFInst_3_n20,
         SubCellInst_LFInst_15_LFInst_3_n19, MCInst_MC0_v1_0_0_,
         MCInst_MC0_v0_2Inst_0_n3, MCInst_MC0_v1_2Inst_0_n3,
         MCInst_MC0_v2_3Inst_0_n6, MCInst_MC0_v2_3Inst_0_n5,
         MCInst_MC0_v3_3Inst_0_n3, MCInst_MC0_v0_2Inst_1_n3,
         MCInst_MC0_v2_1Inst_1_n3, MCInst_MC0_v2_2Inst_1_n6,
         MCInst_MC0_v2_2Inst_1_n5, MCInst_MC0_v3_3Inst_1_n3,
         MCInst_MC0_v1_1Inst_2_n3, MCInst_MC0_v1_2Inst_2_n3,
         MCInst_MC0_v2_1Inst_2_n3, MCInst_MC0_v2_2Inst_2_n3,
         MCInst_MC0_v3_1Inst_2_n3, MCInst_MC0_v1_2Inst_3_n6,
         MCInst_MC0_v1_2Inst_3_n5, MCInst_MC0_v2_2Inst_3_n3,
         MCInst_MC0_v2_3Inst_3_n3, MCInst_MC0_r0Inst_XORInst_0_0_n8,
         MCInst_MC0_r0Inst_XORInst_0_0_n7, MCInst_MC0_r0Inst_XORInst_0_1_n8,
         MCInst_MC0_r0Inst_XORInst_0_1_n7, MCInst_MC0_r0Inst_XORInst_0_2_n8,
         MCInst_MC0_r0Inst_XORInst_0_2_n7, MCInst_MC0_r0Inst_XORInst_0_3_n8,
         MCInst_MC0_r0Inst_XORInst_0_3_n7, MCInst_MC0_r1Inst_XORInst_0_0_n8,
         MCInst_MC0_r1Inst_XORInst_0_0_n7, MCInst_MC0_r1Inst_XORInst_0_1_n8,
         MCInst_MC0_r1Inst_XORInst_0_1_n7, MCInst_MC0_r1Inst_XORInst_0_2_n8,
         MCInst_MC0_r1Inst_XORInst_0_2_n7, MCInst_MC0_r1Inst_XORInst_0_3_n8,
         MCInst_MC0_r1Inst_XORInst_0_3_n7, MCInst_MC0_r2Inst_XORInst_0_0_n8,
         MCInst_MC0_r2Inst_XORInst_0_0_n7, MCInst_MC0_r2Inst_XORInst_0_1_n8,
         MCInst_MC0_r2Inst_XORInst_0_1_n7, MCInst_MC0_r2Inst_XORInst_0_2_n8,
         MCInst_MC0_r2Inst_XORInst_0_2_n7, MCInst_MC0_r2Inst_XORInst_0_3_n8,
         MCInst_MC0_r2Inst_XORInst_0_3_n7, MCInst_MC0_r3Inst_XORInst_0_0_n8,
         MCInst_MC0_r3Inst_XORInst_0_0_n7, MCInst_MC0_r3Inst_XORInst_0_1_n8,
         MCInst_MC0_r3Inst_XORInst_0_1_n7, MCInst_MC0_r3Inst_XORInst_0_2_n8,
         MCInst_MC0_r3Inst_XORInst_0_2_n7, MCInst_MC0_r3Inst_XORInst_0_3_n8,
         MCInst_MC0_r3Inst_XORInst_0_3_n7, MCInst_MC1_v1_0_0_,
         MCInst_MC1_v0_2Inst_0_n3, MCInst_MC1_v1_2Inst_0_n3,
         MCInst_MC1_v2_3Inst_0_n6, MCInst_MC1_v2_3Inst_0_n5,
         MCInst_MC1_v3_3Inst_0_n3, MCInst_MC1_v0_2Inst_1_n3,
         MCInst_MC1_v2_1Inst_1_n3, MCInst_MC1_v2_2Inst_1_n6,
         MCInst_MC1_v2_2Inst_1_n5, MCInst_MC1_v3_3Inst_1_n3,
         MCInst_MC1_v1_1Inst_2_n3, MCInst_MC1_v1_2Inst_2_n3,
         MCInst_MC1_v2_1Inst_2_n3, MCInst_MC1_v2_2Inst_2_n3,
         MCInst_MC1_v3_1Inst_2_n3, MCInst_MC1_v1_2Inst_3_n6,
         MCInst_MC1_v1_2Inst_3_n5, MCInst_MC1_v2_2Inst_3_n3,
         MCInst_MC1_v2_3Inst_3_n3, MCInst_MC1_r0Inst_XORInst_0_0_n8,
         MCInst_MC1_r0Inst_XORInst_0_0_n7, MCInst_MC1_r0Inst_XORInst_0_1_n8,
         MCInst_MC1_r0Inst_XORInst_0_1_n7, MCInst_MC1_r0Inst_XORInst_0_2_n8,
         MCInst_MC1_r0Inst_XORInst_0_2_n7, MCInst_MC1_r0Inst_XORInst_0_3_n8,
         MCInst_MC1_r0Inst_XORInst_0_3_n7, MCInst_MC1_r1Inst_XORInst_0_0_n8,
         MCInst_MC1_r1Inst_XORInst_0_0_n7, MCInst_MC1_r1Inst_XORInst_0_1_n8,
         MCInst_MC1_r1Inst_XORInst_0_1_n7, MCInst_MC1_r1Inst_XORInst_0_2_n8,
         MCInst_MC1_r1Inst_XORInst_0_2_n7, MCInst_MC1_r1Inst_XORInst_0_3_n8,
         MCInst_MC1_r1Inst_XORInst_0_3_n7, MCInst_MC1_r2Inst_XORInst_0_0_n8,
         MCInst_MC1_r2Inst_XORInst_0_0_n7, MCInst_MC1_r2Inst_XORInst_0_1_n8,
         MCInst_MC1_r2Inst_XORInst_0_1_n7, MCInst_MC1_r2Inst_XORInst_0_2_n8,
         MCInst_MC1_r2Inst_XORInst_0_2_n7, MCInst_MC1_r2Inst_XORInst_0_3_n8,
         MCInst_MC1_r2Inst_XORInst_0_3_n7, MCInst_MC1_r3Inst_XORInst_0_0_n8,
         MCInst_MC1_r3Inst_XORInst_0_0_n7, MCInst_MC1_r3Inst_XORInst_0_1_n8,
         MCInst_MC1_r3Inst_XORInst_0_1_n7, MCInst_MC1_r3Inst_XORInst_0_2_n8,
         MCInst_MC1_r3Inst_XORInst_0_2_n7, MCInst_MC1_r3Inst_XORInst_0_3_n8,
         MCInst_MC1_r3Inst_XORInst_0_3_n7, MCInst_MC2_v1_0_0_,
         MCInst_MC2_v0_2Inst_0_n3, MCInst_MC2_v1_2Inst_0_n3,
         MCInst_MC2_v2_3Inst_0_n6, MCInst_MC2_v2_3Inst_0_n5,
         MCInst_MC2_v3_3Inst_0_n3, MCInst_MC2_v0_2Inst_1_n3,
         MCInst_MC2_v2_1Inst_1_n3, MCInst_MC2_v2_2Inst_1_n6,
         MCInst_MC2_v2_2Inst_1_n5, MCInst_MC2_v3_3Inst_1_n3,
         MCInst_MC2_v1_1Inst_2_n3, MCInst_MC2_v1_2Inst_2_n3,
         MCInst_MC2_v2_1Inst_2_n3, MCInst_MC2_v2_2Inst_2_n3,
         MCInst_MC2_v3_1Inst_2_n3, MCInst_MC2_v1_2Inst_3_n6,
         MCInst_MC2_v1_2Inst_3_n5, MCInst_MC2_v2_2Inst_3_n3,
         MCInst_MC2_v2_3Inst_3_n3, MCInst_MC2_r0Inst_XORInst_0_0_n8,
         MCInst_MC2_r0Inst_XORInst_0_0_n7, MCInst_MC2_r0Inst_XORInst_0_1_n8,
         MCInst_MC2_r0Inst_XORInst_0_1_n7, MCInst_MC2_r0Inst_XORInst_0_2_n8,
         MCInst_MC2_r0Inst_XORInst_0_2_n7, MCInst_MC2_r0Inst_XORInst_0_3_n8,
         MCInst_MC2_r0Inst_XORInst_0_3_n7, MCInst_MC2_r1Inst_XORInst_0_0_n8,
         MCInst_MC2_r1Inst_XORInst_0_0_n7, MCInst_MC2_r1Inst_XORInst_0_1_n8,
         MCInst_MC2_r1Inst_XORInst_0_1_n7, MCInst_MC2_r1Inst_XORInst_0_2_n8,
         MCInst_MC2_r1Inst_XORInst_0_2_n7, MCInst_MC2_r1Inst_XORInst_0_3_n8,
         MCInst_MC2_r1Inst_XORInst_0_3_n7, MCInst_MC2_r2Inst_XORInst_0_0_n8,
         MCInst_MC2_r2Inst_XORInst_0_0_n7, MCInst_MC2_r2Inst_XORInst_0_1_n8,
         MCInst_MC2_r2Inst_XORInst_0_1_n7, MCInst_MC2_r2Inst_XORInst_0_2_n8,
         MCInst_MC2_r2Inst_XORInst_0_2_n7, MCInst_MC2_r2Inst_XORInst_0_3_n8,
         MCInst_MC2_r2Inst_XORInst_0_3_n7, MCInst_MC2_r3Inst_XORInst_0_0_n8,
         MCInst_MC2_r3Inst_XORInst_0_0_n7, MCInst_MC2_r3Inst_XORInst_0_1_n8,
         MCInst_MC2_r3Inst_XORInst_0_1_n7, MCInst_MC2_r3Inst_XORInst_0_2_n8,
         MCInst_MC2_r3Inst_XORInst_0_2_n7, MCInst_MC2_r3Inst_XORInst_0_3_n8,
         MCInst_MC2_r3Inst_XORInst_0_3_n7, MCInst_MC3_v1_0_0_,
         MCInst_MC3_v0_2Inst_0_n3, MCInst_MC3_v1_2Inst_0_n3,
         MCInst_MC3_v2_3Inst_0_n6, MCInst_MC3_v2_3Inst_0_n5,
         MCInst_MC3_v3_3Inst_0_n3, MCInst_MC3_v0_2Inst_1_n3,
         MCInst_MC3_v2_1Inst_1_n3, MCInst_MC3_v2_2Inst_1_n6,
         MCInst_MC3_v2_2Inst_1_n5, MCInst_MC3_v3_3Inst_1_n3,
         MCInst_MC3_v1_1Inst_2_n3, MCInst_MC3_v1_2Inst_2_n3,
         MCInst_MC3_v2_1Inst_2_n3, MCInst_MC3_v2_2Inst_2_n3,
         MCInst_MC3_v3_1Inst_2_n3, MCInst_MC3_v1_2Inst_3_n6,
         MCInst_MC3_v1_2Inst_3_n5, MCInst_MC3_v2_2Inst_3_n3,
         MCInst_MC3_v2_3Inst_3_n3, MCInst_MC3_r0Inst_XORInst_0_0_n8,
         MCInst_MC3_r0Inst_XORInst_0_0_n7, MCInst_MC3_r0Inst_XORInst_0_1_n8,
         MCInst_MC3_r0Inst_XORInst_0_1_n7, MCInst_MC3_r0Inst_XORInst_0_2_n8,
         MCInst_MC3_r0Inst_XORInst_0_2_n7, MCInst_MC3_r0Inst_XORInst_0_3_n8,
         MCInst_MC3_r0Inst_XORInst_0_3_n7, MCInst_MC3_r1Inst_XORInst_0_0_n8,
         MCInst_MC3_r1Inst_XORInst_0_0_n7, MCInst_MC3_r1Inst_XORInst_0_1_n8,
         MCInst_MC3_r1Inst_XORInst_0_1_n7, MCInst_MC3_r1Inst_XORInst_0_2_n8,
         MCInst_MC3_r1Inst_XORInst_0_2_n7, MCInst_MC3_r1Inst_XORInst_0_3_n8,
         MCInst_MC3_r1Inst_XORInst_0_3_n7, MCInst_MC3_r2Inst_XORInst_0_0_n8,
         MCInst_MC3_r2Inst_XORInst_0_0_n7, MCInst_MC3_r2Inst_XORInst_0_1_n8,
         MCInst_MC3_r2Inst_XORInst_0_1_n7, MCInst_MC3_r2Inst_XORInst_0_2_n8,
         MCInst_MC3_r2Inst_XORInst_0_2_n7, MCInst_MC3_r2Inst_XORInst_0_3_n8,
         MCInst_MC3_r2Inst_XORInst_0_3_n7, MCInst_MC3_r3Inst_XORInst_0_0_n8,
         MCInst_MC3_r3Inst_XORInst_0_0_n7, MCInst_MC3_r3Inst_XORInst_0_1_n8,
         MCInst_MC3_r3Inst_XORInst_0_1_n7, MCInst_MC3_r3Inst_XORInst_0_2_n8,
         MCInst_MC3_r3Inst_XORInst_0_2_n7, MCInst_MC3_r3Inst_XORInst_0_3_n8,
         MCInst_MC3_r3Inst_XORInst_0_3_n7, SubCellInst2_LFInst_0_LFInst_0_n7,
         SubCellInst2_LFInst_0_LFInst_0_n6, SubCellInst2_LFInst_0_LFInst_0_n5,
         SubCellInst2_LFInst_0_LFInst_0_n8, SubCellInst2_LFInst_0_LFInst_1_n26,
         SubCellInst2_LFInst_0_LFInst_1_n25,
         SubCellInst2_LFInst_0_LFInst_1_n24,
         SubCellInst2_LFInst_0_LFInst_1_n23,
         SubCellInst2_LFInst_0_LFInst_1_n22,
         SubCellInst2_LFInst_0_LFInst_1_n21,
         SubCellInst2_LFInst_0_LFInst_1_n20,
         SubCellInst2_LFInst_0_LFInst_1_n19,
         SubCellInst2_LFInst_0_LFInst_1_n18,
         SubCellInst2_LFInst_0_LFInst_2_n28,
         SubCellInst2_LFInst_0_LFInst_2_n27,
         SubCellInst2_LFInst_0_LFInst_2_n26,
         SubCellInst2_LFInst_0_LFInst_2_n25,
         SubCellInst2_LFInst_0_LFInst_2_n24,
         SubCellInst2_LFInst_0_LFInst_2_n23,
         SubCellInst2_LFInst_0_LFInst_2_n22,
         SubCellInst2_LFInst_0_LFInst_3_n26,
         SubCellInst2_LFInst_0_LFInst_3_n25,
         SubCellInst2_LFInst_0_LFInst_3_n24,
         SubCellInst2_LFInst_0_LFInst_3_n23,
         SubCellInst2_LFInst_0_LFInst_3_n22,
         SubCellInst2_LFInst_0_LFInst_3_n21,
         SubCellInst2_LFInst_0_LFInst_3_n20,
         SubCellInst2_LFInst_0_LFInst_3_n19, SubCellInst2_LFInst_1_LFInst_0_n7,
         SubCellInst2_LFInst_1_LFInst_0_n6, SubCellInst2_LFInst_1_LFInst_0_n5,
         SubCellInst2_LFInst_1_LFInst_0_n8, SubCellInst2_LFInst_1_LFInst_1_n26,
         SubCellInst2_LFInst_1_LFInst_1_n25,
         SubCellInst2_LFInst_1_LFInst_1_n24,
         SubCellInst2_LFInst_1_LFInst_1_n23,
         SubCellInst2_LFInst_1_LFInst_1_n22,
         SubCellInst2_LFInst_1_LFInst_1_n21,
         SubCellInst2_LFInst_1_LFInst_1_n20,
         SubCellInst2_LFInst_1_LFInst_1_n19,
         SubCellInst2_LFInst_1_LFInst_1_n18,
         SubCellInst2_LFInst_1_LFInst_2_n29,
         SubCellInst2_LFInst_1_LFInst_2_n28,
         SubCellInst2_LFInst_1_LFInst_2_n27,
         SubCellInst2_LFInst_1_LFInst_2_n26,
         SubCellInst2_LFInst_1_LFInst_2_n25,
         SubCellInst2_LFInst_1_LFInst_2_n24,
         SubCellInst2_LFInst_1_LFInst_2_n23,
         SubCellInst2_LFInst_1_LFInst_2_n22,
         SubCellInst2_LFInst_1_LFInst_3_n26,
         SubCellInst2_LFInst_1_LFInst_3_n25,
         SubCellInst2_LFInst_1_LFInst_3_n24,
         SubCellInst2_LFInst_1_LFInst_3_n23,
         SubCellInst2_LFInst_1_LFInst_3_n22,
         SubCellInst2_LFInst_1_LFInst_3_n21,
         SubCellInst2_LFInst_1_LFInst_3_n20,
         SubCellInst2_LFInst_1_LFInst_3_n19, SubCellInst2_LFInst_2_LFInst_0_n7,
         SubCellInst2_LFInst_2_LFInst_0_n6, SubCellInst2_LFInst_2_LFInst_0_n5,
         SubCellInst2_LFInst_2_LFInst_0_n8, SubCellInst2_LFInst_2_LFInst_1_n26,
         SubCellInst2_LFInst_2_LFInst_1_n25,
         SubCellInst2_LFInst_2_LFInst_1_n24,
         SubCellInst2_LFInst_2_LFInst_1_n23,
         SubCellInst2_LFInst_2_LFInst_1_n22,
         SubCellInst2_LFInst_2_LFInst_1_n21,
         SubCellInst2_LFInst_2_LFInst_1_n20,
         SubCellInst2_LFInst_2_LFInst_1_n19,
         SubCellInst2_LFInst_2_LFInst_1_n18,
         SubCellInst2_LFInst_2_LFInst_2_n28,
         SubCellInst2_LFInst_2_LFInst_2_n27,
         SubCellInst2_LFInst_2_LFInst_2_n26,
         SubCellInst2_LFInst_2_LFInst_2_n25,
         SubCellInst2_LFInst_2_LFInst_2_n24,
         SubCellInst2_LFInst_2_LFInst_2_n23,
         SubCellInst2_LFInst_2_LFInst_2_n22,
         SubCellInst2_LFInst_2_LFInst_3_n26,
         SubCellInst2_LFInst_2_LFInst_3_n25,
         SubCellInst2_LFInst_2_LFInst_3_n24,
         SubCellInst2_LFInst_2_LFInst_3_n23,
         SubCellInst2_LFInst_2_LFInst_3_n22,
         SubCellInst2_LFInst_2_LFInst_3_n21,
         SubCellInst2_LFInst_2_LFInst_3_n20,
         SubCellInst2_LFInst_2_LFInst_3_n19, SubCellInst2_LFInst_3_LFInst_0_n7,
         SubCellInst2_LFInst_3_LFInst_0_n6, SubCellInst2_LFInst_3_LFInst_0_n5,
         SubCellInst2_LFInst_3_LFInst_0_n8, SubCellInst2_LFInst_3_LFInst_1_n26,
         SubCellInst2_LFInst_3_LFInst_1_n25,
         SubCellInst2_LFInst_3_LFInst_1_n24,
         SubCellInst2_LFInst_3_LFInst_1_n23,
         SubCellInst2_LFInst_3_LFInst_1_n22,
         SubCellInst2_LFInst_3_LFInst_1_n21,
         SubCellInst2_LFInst_3_LFInst_1_n20,
         SubCellInst2_LFInst_3_LFInst_1_n19,
         SubCellInst2_LFInst_3_LFInst_1_n18,
         SubCellInst2_LFInst_3_LFInst_2_n28,
         SubCellInst2_LFInst_3_LFInst_2_n27,
         SubCellInst2_LFInst_3_LFInst_2_n26,
         SubCellInst2_LFInst_3_LFInst_2_n25,
         SubCellInst2_LFInst_3_LFInst_2_n24,
         SubCellInst2_LFInst_3_LFInst_2_n23,
         SubCellInst2_LFInst_3_LFInst_2_n22,
         SubCellInst2_LFInst_3_LFInst_3_n26,
         SubCellInst2_LFInst_3_LFInst_3_n25,
         SubCellInst2_LFInst_3_LFInst_3_n24,
         SubCellInst2_LFInst_3_LFInst_3_n23,
         SubCellInst2_LFInst_3_LFInst_3_n22,
         SubCellInst2_LFInst_3_LFInst_3_n21,
         SubCellInst2_LFInst_3_LFInst_3_n20,
         SubCellInst2_LFInst_3_LFInst_3_n19, SubCellInst2_LFInst_4_LFInst_0_n6,
         SubCellInst2_LFInst_4_LFInst_0_n5, SubCellInst2_LFInst_4_LFInst_0_n4,
         SubCellInst2_LFInst_4_LFInst_1_n26,
         SubCellInst2_LFInst_4_LFInst_1_n25,
         SubCellInst2_LFInst_4_LFInst_1_n24,
         SubCellInst2_LFInst_4_LFInst_1_n23,
         SubCellInst2_LFInst_4_LFInst_1_n22,
         SubCellInst2_LFInst_4_LFInst_1_n21,
         SubCellInst2_LFInst_4_LFInst_1_n20,
         SubCellInst2_LFInst_4_LFInst_1_n19,
         SubCellInst2_LFInst_4_LFInst_1_n18,
         SubCellInst2_LFInst_4_LFInst_2_n29,
         SubCellInst2_LFInst_4_LFInst_2_n28,
         SubCellInst2_LFInst_4_LFInst_2_n27,
         SubCellInst2_LFInst_4_LFInst_2_n26,
         SubCellInst2_LFInst_4_LFInst_2_n25,
         SubCellInst2_LFInst_4_LFInst_2_n24,
         SubCellInst2_LFInst_4_LFInst_2_n23,
         SubCellInst2_LFInst_4_LFInst_2_n22,
         SubCellInst2_LFInst_4_LFInst_3_n26,
         SubCellInst2_LFInst_4_LFInst_3_n25,
         SubCellInst2_LFInst_4_LFInst_3_n24,
         SubCellInst2_LFInst_4_LFInst_3_n23,
         SubCellInst2_LFInst_4_LFInst_3_n22,
         SubCellInst2_LFInst_4_LFInst_3_n21,
         SubCellInst2_LFInst_4_LFInst_3_n20,
         SubCellInst2_LFInst_4_LFInst_3_n19, SubCellInst2_LFInst_5_LFInst_0_n6,
         SubCellInst2_LFInst_5_LFInst_0_n5, SubCellInst2_LFInst_5_LFInst_0_n4,
         SubCellInst2_LFInst_5_LFInst_1_n26,
         SubCellInst2_LFInst_5_LFInst_1_n25,
         SubCellInst2_LFInst_5_LFInst_1_n24,
         SubCellInst2_LFInst_5_LFInst_1_n23,
         SubCellInst2_LFInst_5_LFInst_1_n22,
         SubCellInst2_LFInst_5_LFInst_1_n21,
         SubCellInst2_LFInst_5_LFInst_1_n20,
         SubCellInst2_LFInst_5_LFInst_1_n19,
         SubCellInst2_LFInst_5_LFInst_1_n18,
         SubCellInst2_LFInst_5_LFInst_2_n29,
         SubCellInst2_LFInst_5_LFInst_2_n28,
         SubCellInst2_LFInst_5_LFInst_2_n27,
         SubCellInst2_LFInst_5_LFInst_2_n26,
         SubCellInst2_LFInst_5_LFInst_2_n25,
         SubCellInst2_LFInst_5_LFInst_2_n24,
         SubCellInst2_LFInst_5_LFInst_2_n23,
         SubCellInst2_LFInst_5_LFInst_2_n22,
         SubCellInst2_LFInst_5_LFInst_3_n26,
         SubCellInst2_LFInst_5_LFInst_3_n25,
         SubCellInst2_LFInst_5_LFInst_3_n24,
         SubCellInst2_LFInst_5_LFInst_3_n23,
         SubCellInst2_LFInst_5_LFInst_3_n22,
         SubCellInst2_LFInst_5_LFInst_3_n21,
         SubCellInst2_LFInst_5_LFInst_3_n20,
         SubCellInst2_LFInst_5_LFInst_3_n19, SubCellInst2_LFInst_6_LFInst_0_n6,
         SubCellInst2_LFInst_6_LFInst_0_n5, SubCellInst2_LFInst_6_LFInst_0_n4,
         SubCellInst2_LFInst_6_LFInst_1_n26,
         SubCellInst2_LFInst_6_LFInst_1_n25,
         SubCellInst2_LFInst_6_LFInst_1_n24,
         SubCellInst2_LFInst_6_LFInst_1_n23,
         SubCellInst2_LFInst_6_LFInst_1_n22,
         SubCellInst2_LFInst_6_LFInst_1_n21,
         SubCellInst2_LFInst_6_LFInst_1_n20,
         SubCellInst2_LFInst_6_LFInst_1_n19,
         SubCellInst2_LFInst_6_LFInst_1_n18,
         SubCellInst2_LFInst_6_LFInst_2_n29,
         SubCellInst2_LFInst_6_LFInst_2_n28,
         SubCellInst2_LFInst_6_LFInst_2_n27,
         SubCellInst2_LFInst_6_LFInst_2_n26,
         SubCellInst2_LFInst_6_LFInst_2_n25,
         SubCellInst2_LFInst_6_LFInst_2_n24,
         SubCellInst2_LFInst_6_LFInst_2_n23,
         SubCellInst2_LFInst_6_LFInst_2_n22,
         SubCellInst2_LFInst_6_LFInst_3_n26,
         SubCellInst2_LFInst_6_LFInst_3_n25,
         SubCellInst2_LFInst_6_LFInst_3_n24,
         SubCellInst2_LFInst_6_LFInst_3_n23,
         SubCellInst2_LFInst_6_LFInst_3_n22,
         SubCellInst2_LFInst_6_LFInst_3_n21,
         SubCellInst2_LFInst_6_LFInst_3_n20,
         SubCellInst2_LFInst_6_LFInst_3_n19, SubCellInst2_LFInst_7_LFInst_0_n6,
         SubCellInst2_LFInst_7_LFInst_0_n5, SubCellInst2_LFInst_7_LFInst_0_n4,
         SubCellInst2_LFInst_7_LFInst_1_n26,
         SubCellInst2_LFInst_7_LFInst_1_n25,
         SubCellInst2_LFInst_7_LFInst_1_n24,
         SubCellInst2_LFInst_7_LFInst_1_n23,
         SubCellInst2_LFInst_7_LFInst_1_n22,
         SubCellInst2_LFInst_7_LFInst_1_n21,
         SubCellInst2_LFInst_7_LFInst_1_n20,
         SubCellInst2_LFInst_7_LFInst_1_n19,
         SubCellInst2_LFInst_7_LFInst_1_n18,
         SubCellInst2_LFInst_7_LFInst_2_n29,
         SubCellInst2_LFInst_7_LFInst_2_n28,
         SubCellInst2_LFInst_7_LFInst_2_n27,
         SubCellInst2_LFInst_7_LFInst_2_n26,
         SubCellInst2_LFInst_7_LFInst_2_n25,
         SubCellInst2_LFInst_7_LFInst_2_n24,
         SubCellInst2_LFInst_7_LFInst_2_n23,
         SubCellInst2_LFInst_7_LFInst_2_n22,
         SubCellInst2_LFInst_7_LFInst_3_n26,
         SubCellInst2_LFInst_7_LFInst_3_n25,
         SubCellInst2_LFInst_7_LFInst_3_n24,
         SubCellInst2_LFInst_7_LFInst_3_n23,
         SubCellInst2_LFInst_7_LFInst_3_n22,
         SubCellInst2_LFInst_7_LFInst_3_n21,
         SubCellInst2_LFInst_7_LFInst_3_n20,
         SubCellInst2_LFInst_7_LFInst_3_n19, SubCellInst2_LFInst_8_LFInst_0_n9,
         SubCellInst2_LFInst_8_LFInst_0_n8, SubCellInst2_LFInst_8_LFInst_0_n7,
         SubCellInst2_LFInst_8_LFInst_0_n10,
         SubCellInst2_LFInst_8_LFInst_1_n26,
         SubCellInst2_LFInst_8_LFInst_1_n25,
         SubCellInst2_LFInst_8_LFInst_1_n24,
         SubCellInst2_LFInst_8_LFInst_1_n23,
         SubCellInst2_LFInst_8_LFInst_1_n22,
         SubCellInst2_LFInst_8_LFInst_1_n21,
         SubCellInst2_LFInst_8_LFInst_1_n20,
         SubCellInst2_LFInst_8_LFInst_1_n19,
         SubCellInst2_LFInst_8_LFInst_1_n18,
         SubCellInst2_LFInst_8_LFInst_2_n29,
         SubCellInst2_LFInst_8_LFInst_2_n28,
         SubCellInst2_LFInst_8_LFInst_2_n27,
         SubCellInst2_LFInst_8_LFInst_2_n26,
         SubCellInst2_LFInst_8_LFInst_2_n25,
         SubCellInst2_LFInst_8_LFInst_2_n24,
         SubCellInst2_LFInst_8_LFInst_2_n23,
         SubCellInst2_LFInst_8_LFInst_2_n22,
         SubCellInst2_LFInst_8_LFInst_3_n26,
         SubCellInst2_LFInst_8_LFInst_3_n25,
         SubCellInst2_LFInst_8_LFInst_3_n24,
         SubCellInst2_LFInst_8_LFInst_3_n23,
         SubCellInst2_LFInst_8_LFInst_3_n22,
         SubCellInst2_LFInst_8_LFInst_3_n21,
         SubCellInst2_LFInst_8_LFInst_3_n20,
         SubCellInst2_LFInst_8_LFInst_3_n19,
         SubCellInst2_LFInst_9_LFInst_0_n10, SubCellInst2_LFInst_9_LFInst_0_n9,
         SubCellInst2_LFInst_9_LFInst_0_n8, SubCellInst2_LFInst_9_LFInst_0_n7,
         SubCellInst2_LFInst_9_LFInst_1_n26,
         SubCellInst2_LFInst_9_LFInst_1_n25,
         SubCellInst2_LFInst_9_LFInst_1_n24,
         SubCellInst2_LFInst_9_LFInst_1_n23,
         SubCellInst2_LFInst_9_LFInst_1_n22,
         SubCellInst2_LFInst_9_LFInst_1_n21,
         SubCellInst2_LFInst_9_LFInst_1_n20,
         SubCellInst2_LFInst_9_LFInst_1_n19,
         SubCellInst2_LFInst_9_LFInst_1_n18,
         SubCellInst2_LFInst_9_LFInst_2_n29,
         SubCellInst2_LFInst_9_LFInst_2_n28,
         SubCellInst2_LFInst_9_LFInst_2_n27,
         SubCellInst2_LFInst_9_LFInst_2_n26,
         SubCellInst2_LFInst_9_LFInst_2_n25,
         SubCellInst2_LFInst_9_LFInst_2_n24,
         SubCellInst2_LFInst_9_LFInst_2_n23,
         SubCellInst2_LFInst_9_LFInst_2_n22,
         SubCellInst2_LFInst_9_LFInst_3_n26,
         SubCellInst2_LFInst_9_LFInst_3_n25,
         SubCellInst2_LFInst_9_LFInst_3_n24,
         SubCellInst2_LFInst_9_LFInst_3_n23,
         SubCellInst2_LFInst_9_LFInst_3_n22,
         SubCellInst2_LFInst_9_LFInst_3_n21,
         SubCellInst2_LFInst_9_LFInst_3_n20,
         SubCellInst2_LFInst_9_LFInst_3_n19,
         SubCellInst2_LFInst_10_LFInst_0_n10,
         SubCellInst2_LFInst_10_LFInst_0_n9,
         SubCellInst2_LFInst_10_LFInst_0_n8,
         SubCellInst2_LFInst_10_LFInst_0_n7,
         SubCellInst2_LFInst_10_LFInst_1_n26,
         SubCellInst2_LFInst_10_LFInst_1_n25,
         SubCellInst2_LFInst_10_LFInst_1_n24,
         SubCellInst2_LFInst_10_LFInst_1_n23,
         SubCellInst2_LFInst_10_LFInst_1_n22,
         SubCellInst2_LFInst_10_LFInst_1_n21,
         SubCellInst2_LFInst_10_LFInst_1_n20,
         SubCellInst2_LFInst_10_LFInst_1_n19,
         SubCellInst2_LFInst_10_LFInst_1_n18,
         SubCellInst2_LFInst_10_LFInst_2_n29,
         SubCellInst2_LFInst_10_LFInst_2_n28,
         SubCellInst2_LFInst_10_LFInst_2_n27,
         SubCellInst2_LFInst_10_LFInst_2_n26,
         SubCellInst2_LFInst_10_LFInst_2_n25,
         SubCellInst2_LFInst_10_LFInst_2_n24,
         SubCellInst2_LFInst_10_LFInst_2_n23,
         SubCellInst2_LFInst_10_LFInst_2_n22,
         SubCellInst2_LFInst_10_LFInst_3_n26,
         SubCellInst2_LFInst_10_LFInst_3_n25,
         SubCellInst2_LFInst_10_LFInst_3_n24,
         SubCellInst2_LFInst_10_LFInst_3_n23,
         SubCellInst2_LFInst_10_LFInst_3_n22,
         SubCellInst2_LFInst_10_LFInst_3_n21,
         SubCellInst2_LFInst_10_LFInst_3_n20,
         SubCellInst2_LFInst_10_LFInst_3_n19,
         SubCellInst2_LFInst_11_LFInst_0_n10,
         SubCellInst2_LFInst_11_LFInst_0_n9,
         SubCellInst2_LFInst_11_LFInst_0_n8,
         SubCellInst2_LFInst_11_LFInst_0_n7,
         SubCellInst2_LFInst_11_LFInst_1_n26,
         SubCellInst2_LFInst_11_LFInst_1_n25,
         SubCellInst2_LFInst_11_LFInst_1_n24,
         SubCellInst2_LFInst_11_LFInst_1_n23,
         SubCellInst2_LFInst_11_LFInst_1_n22,
         SubCellInst2_LFInst_11_LFInst_1_n21,
         SubCellInst2_LFInst_11_LFInst_1_n20,
         SubCellInst2_LFInst_11_LFInst_1_n19,
         SubCellInst2_LFInst_11_LFInst_1_n18,
         SubCellInst2_LFInst_11_LFInst_2_n28,
         SubCellInst2_LFInst_11_LFInst_2_n27,
         SubCellInst2_LFInst_11_LFInst_2_n26,
         SubCellInst2_LFInst_11_LFInst_2_n25,
         SubCellInst2_LFInst_11_LFInst_2_n24,
         SubCellInst2_LFInst_11_LFInst_2_n23,
         SubCellInst2_LFInst_11_LFInst_2_n22,
         SubCellInst2_LFInst_11_LFInst_3_n26,
         SubCellInst2_LFInst_11_LFInst_3_n25,
         SubCellInst2_LFInst_11_LFInst_3_n24,
         SubCellInst2_LFInst_11_LFInst_3_n23,
         SubCellInst2_LFInst_11_LFInst_3_n22,
         SubCellInst2_LFInst_11_LFInst_3_n21,
         SubCellInst2_LFInst_11_LFInst_3_n20,
         SubCellInst2_LFInst_11_LFInst_3_n19,
         SubCellInst2_LFInst_12_LFInst_0_n7,
         SubCellInst2_LFInst_12_LFInst_0_n6,
         SubCellInst2_LFInst_12_LFInst_0_n5,
         SubCellInst2_LFInst_12_LFInst_0_n8,
         SubCellInst2_LFInst_12_LFInst_1_n26,
         SubCellInst2_LFInst_12_LFInst_1_n25,
         SubCellInst2_LFInst_12_LFInst_1_n24,
         SubCellInst2_LFInst_12_LFInst_1_n23,
         SubCellInst2_LFInst_12_LFInst_1_n22,
         SubCellInst2_LFInst_12_LFInst_1_n21,
         SubCellInst2_LFInst_12_LFInst_1_n20,
         SubCellInst2_LFInst_12_LFInst_1_n19,
         SubCellInst2_LFInst_12_LFInst_1_n18,
         SubCellInst2_LFInst_12_LFInst_2_n29,
         SubCellInst2_LFInst_12_LFInst_2_n28,
         SubCellInst2_LFInst_12_LFInst_2_n27,
         SubCellInst2_LFInst_12_LFInst_2_n26,
         SubCellInst2_LFInst_12_LFInst_2_n25,
         SubCellInst2_LFInst_12_LFInst_2_n24,
         SubCellInst2_LFInst_12_LFInst_2_n23,
         SubCellInst2_LFInst_12_LFInst_2_n22,
         SubCellInst2_LFInst_12_LFInst_3_n26,
         SubCellInst2_LFInst_12_LFInst_3_n25,
         SubCellInst2_LFInst_12_LFInst_3_n24,
         SubCellInst2_LFInst_12_LFInst_3_n23,
         SubCellInst2_LFInst_12_LFInst_3_n22,
         SubCellInst2_LFInst_12_LFInst_3_n21,
         SubCellInst2_LFInst_12_LFInst_3_n20,
         SubCellInst2_LFInst_12_LFInst_3_n19,
         SubCellInst2_LFInst_13_LFInst_0_n7,
         SubCellInst2_LFInst_13_LFInst_0_n6,
         SubCellInst2_LFInst_13_LFInst_0_n5,
         SubCellInst2_LFInst_13_LFInst_0_n8,
         SubCellInst2_LFInst_13_LFInst_1_n26,
         SubCellInst2_LFInst_13_LFInst_1_n25,
         SubCellInst2_LFInst_13_LFInst_1_n24,
         SubCellInst2_LFInst_13_LFInst_1_n23,
         SubCellInst2_LFInst_13_LFInst_1_n22,
         SubCellInst2_LFInst_13_LFInst_1_n21,
         SubCellInst2_LFInst_13_LFInst_1_n20,
         SubCellInst2_LFInst_13_LFInst_1_n19,
         SubCellInst2_LFInst_13_LFInst_1_n18,
         SubCellInst2_LFInst_13_LFInst_2_n29,
         SubCellInst2_LFInst_13_LFInst_2_n28,
         SubCellInst2_LFInst_13_LFInst_2_n27,
         SubCellInst2_LFInst_13_LFInst_2_n26,
         SubCellInst2_LFInst_13_LFInst_2_n25,
         SubCellInst2_LFInst_13_LFInst_2_n24,
         SubCellInst2_LFInst_13_LFInst_2_n23,
         SubCellInst2_LFInst_13_LFInst_2_n22,
         SubCellInst2_LFInst_13_LFInst_3_n26,
         SubCellInst2_LFInst_13_LFInst_3_n25,
         SubCellInst2_LFInst_13_LFInst_3_n24,
         SubCellInst2_LFInst_13_LFInst_3_n23,
         SubCellInst2_LFInst_13_LFInst_3_n22,
         SubCellInst2_LFInst_13_LFInst_3_n21,
         SubCellInst2_LFInst_13_LFInst_3_n20,
         SubCellInst2_LFInst_13_LFInst_3_n19,
         SubCellInst2_LFInst_14_LFInst_0_n7,
         SubCellInst2_LFInst_14_LFInst_0_n6,
         SubCellInst2_LFInst_14_LFInst_0_n5,
         SubCellInst2_LFInst_14_LFInst_0_n8,
         SubCellInst2_LFInst_14_LFInst_1_n26,
         SubCellInst2_LFInst_14_LFInst_1_n25,
         SubCellInst2_LFInst_14_LFInst_1_n24,
         SubCellInst2_LFInst_14_LFInst_1_n23,
         SubCellInst2_LFInst_14_LFInst_1_n22,
         SubCellInst2_LFInst_14_LFInst_1_n21,
         SubCellInst2_LFInst_14_LFInst_1_n20,
         SubCellInst2_LFInst_14_LFInst_1_n19,
         SubCellInst2_LFInst_14_LFInst_1_n18,
         SubCellInst2_LFInst_14_LFInst_2_n29,
         SubCellInst2_LFInst_14_LFInst_2_n28,
         SubCellInst2_LFInst_14_LFInst_2_n27,
         SubCellInst2_LFInst_14_LFInst_2_n26,
         SubCellInst2_LFInst_14_LFInst_2_n25,
         SubCellInst2_LFInst_14_LFInst_2_n24,
         SubCellInst2_LFInst_14_LFInst_2_n23,
         SubCellInst2_LFInst_14_LFInst_2_n22,
         SubCellInst2_LFInst_14_LFInst_3_n26,
         SubCellInst2_LFInst_14_LFInst_3_n25,
         SubCellInst2_LFInst_14_LFInst_3_n24,
         SubCellInst2_LFInst_14_LFInst_3_n23,
         SubCellInst2_LFInst_14_LFInst_3_n22,
         SubCellInst2_LFInst_14_LFInst_3_n21,
         SubCellInst2_LFInst_14_LFInst_3_n20,
         SubCellInst2_LFInst_14_LFInst_3_n19,
         SubCellInst2_LFInst_15_LFInst_0_n7,
         SubCellInst2_LFInst_15_LFInst_0_n6,
         SubCellInst2_LFInst_15_LFInst_0_n5,
         SubCellInst2_LFInst_15_LFInst_0_n8,
         SubCellInst2_LFInst_15_LFInst_1_n26,
         SubCellInst2_LFInst_15_LFInst_1_n25,
         SubCellInst2_LFInst_15_LFInst_1_n24,
         SubCellInst2_LFInst_15_LFInst_1_n23,
         SubCellInst2_LFInst_15_LFInst_1_n22,
         SubCellInst2_LFInst_15_LFInst_1_n21,
         SubCellInst2_LFInst_15_LFInst_1_n20,
         SubCellInst2_LFInst_15_LFInst_1_n19,
         SubCellInst2_LFInst_15_LFInst_1_n18,
         SubCellInst2_LFInst_15_LFInst_2_n29,
         SubCellInst2_LFInst_15_LFInst_2_n28,
         SubCellInst2_LFInst_15_LFInst_2_n27,
         SubCellInst2_LFInst_15_LFInst_2_n26,
         SubCellInst2_LFInst_15_LFInst_2_n25,
         SubCellInst2_LFInst_15_LFInst_2_n24,
         SubCellInst2_LFInst_15_LFInst_2_n23,
         SubCellInst2_LFInst_15_LFInst_2_n22,
         SubCellInst2_LFInst_15_LFInst_3_n26,
         SubCellInst2_LFInst_15_LFInst_3_n25,
         SubCellInst2_LFInst_15_LFInst_3_n24,
         SubCellInst2_LFInst_15_LFInst_3_n23,
         SubCellInst2_LFInst_15_LFInst_3_n22,
         SubCellInst2_LFInst_15_LFInst_3_n21,
         SubCellInst2_LFInst_15_LFInst_3_n20,
         SubCellInst2_LFInst_15_LFInst_3_n19, MCInst2_MC0_v1_0_0_,
         MCInst2_MC0_v0_2Inst_0_n3, MCInst2_MC0_v1_2Inst_0_n3,
         MCInst2_MC0_v2_3Inst_0_n6, MCInst2_MC0_v2_3Inst_0_n5,
         MCInst2_MC0_v3_3Inst_0_n3, MCInst2_MC0_v0_2Inst_1_n3,
         MCInst2_MC0_v2_1Inst_1_n3, MCInst2_MC0_v2_2Inst_1_n6,
         MCInst2_MC0_v2_2Inst_1_n5, MCInst2_MC0_v3_3Inst_1_n3,
         MCInst2_MC0_v1_1Inst_2_n3, MCInst2_MC0_v1_2Inst_2_n3,
         MCInst2_MC0_v2_1Inst_2_n3, MCInst2_MC0_v2_2Inst_2_n3,
         MCInst2_MC0_v3_1Inst_2_n3, MCInst2_MC0_v1_2Inst_3_n6,
         MCInst2_MC0_v1_2Inst_3_n5, MCInst2_MC0_v2_2Inst_3_n3,
         MCInst2_MC0_v2_3Inst_3_n3, MCInst2_MC0_r0Inst_XORInst_0_0_n8,
         MCInst2_MC0_r0Inst_XORInst_0_0_n7, MCInst2_MC0_r0Inst_XORInst_0_1_n8,
         MCInst2_MC0_r0Inst_XORInst_0_1_n7, MCInst2_MC0_r0Inst_XORInst_0_2_n8,
         MCInst2_MC0_r0Inst_XORInst_0_2_n7, MCInst2_MC0_r0Inst_XORInst_0_3_n8,
         MCInst2_MC0_r0Inst_XORInst_0_3_n7, MCInst2_MC0_r1Inst_XORInst_0_0_n8,
         MCInst2_MC0_r1Inst_XORInst_0_0_n7, MCInst2_MC0_r1Inst_XORInst_0_1_n8,
         MCInst2_MC0_r1Inst_XORInst_0_1_n7, MCInst2_MC0_r1Inst_XORInst_0_2_n8,
         MCInst2_MC0_r1Inst_XORInst_0_2_n7, MCInst2_MC0_r1Inst_XORInst_0_3_n8,
         MCInst2_MC0_r1Inst_XORInst_0_3_n7, MCInst2_MC0_r2Inst_XORInst_0_0_n8,
         MCInst2_MC0_r2Inst_XORInst_0_0_n7, MCInst2_MC0_r2Inst_XORInst_0_1_n8,
         MCInst2_MC0_r2Inst_XORInst_0_1_n7, MCInst2_MC0_r2Inst_XORInst_0_2_n8,
         MCInst2_MC0_r2Inst_XORInst_0_2_n7, MCInst2_MC0_r2Inst_XORInst_0_3_n8,
         MCInst2_MC0_r2Inst_XORInst_0_3_n7, MCInst2_MC0_r3Inst_XORInst_0_0_n8,
         MCInst2_MC0_r3Inst_XORInst_0_0_n7, MCInst2_MC0_r3Inst_XORInst_0_1_n8,
         MCInst2_MC0_r3Inst_XORInst_0_1_n7, MCInst2_MC0_r3Inst_XORInst_0_2_n8,
         MCInst2_MC0_r3Inst_XORInst_0_2_n7, MCInst2_MC0_r3Inst_XORInst_0_3_n8,
         MCInst2_MC0_r3Inst_XORInst_0_3_n7, MCInst2_MC1_v1_0_0_,
         MCInst2_MC1_v0_2Inst_0_n3, MCInst2_MC1_v1_2Inst_0_n3,
         MCInst2_MC1_v2_3Inst_0_n6, MCInst2_MC1_v2_3Inst_0_n5,
         MCInst2_MC1_v3_3Inst_0_n3, MCInst2_MC1_v0_2Inst_1_n3,
         MCInst2_MC1_v2_1Inst_1_n3, MCInst2_MC1_v2_2Inst_1_n6,
         MCInst2_MC1_v2_2Inst_1_n5, MCInst2_MC1_v3_3Inst_1_n3,
         MCInst2_MC1_v1_1Inst_2_n3, MCInst2_MC1_v1_2Inst_2_n3,
         MCInst2_MC1_v2_1Inst_2_n3, MCInst2_MC1_v2_2Inst_2_n3,
         MCInst2_MC1_v3_1Inst_2_n3, MCInst2_MC1_v1_2Inst_3_n6,
         MCInst2_MC1_v1_2Inst_3_n5, MCInst2_MC1_v2_2Inst_3_n3,
         MCInst2_MC1_v2_3Inst_3_n3, MCInst2_MC1_r0Inst_XORInst_0_0_n8,
         MCInst2_MC1_r0Inst_XORInst_0_0_n7, MCInst2_MC1_r0Inst_XORInst_0_1_n8,
         MCInst2_MC1_r0Inst_XORInst_0_1_n7, MCInst2_MC1_r0Inst_XORInst_0_2_n8,
         MCInst2_MC1_r0Inst_XORInst_0_2_n7, MCInst2_MC1_r0Inst_XORInst_0_3_n8,
         MCInst2_MC1_r0Inst_XORInst_0_3_n7, MCInst2_MC1_r1Inst_XORInst_0_0_n8,
         MCInst2_MC1_r1Inst_XORInst_0_0_n7, MCInst2_MC1_r1Inst_XORInst_0_1_n8,
         MCInst2_MC1_r1Inst_XORInst_0_1_n7, MCInst2_MC1_r1Inst_XORInst_0_2_n8,
         MCInst2_MC1_r1Inst_XORInst_0_2_n7, MCInst2_MC1_r1Inst_XORInst_0_3_n8,
         MCInst2_MC1_r1Inst_XORInst_0_3_n7, MCInst2_MC1_r2Inst_XORInst_0_0_n8,
         MCInst2_MC1_r2Inst_XORInst_0_0_n7, MCInst2_MC1_r2Inst_XORInst_0_1_n8,
         MCInst2_MC1_r2Inst_XORInst_0_1_n7, MCInst2_MC1_r2Inst_XORInst_0_2_n8,
         MCInst2_MC1_r2Inst_XORInst_0_2_n7, MCInst2_MC1_r2Inst_XORInst_0_3_n8,
         MCInst2_MC1_r2Inst_XORInst_0_3_n7, MCInst2_MC1_r3Inst_XORInst_0_0_n8,
         MCInst2_MC1_r3Inst_XORInst_0_0_n7, MCInst2_MC1_r3Inst_XORInst_0_1_n8,
         MCInst2_MC1_r3Inst_XORInst_0_1_n7, MCInst2_MC1_r3Inst_XORInst_0_2_n8,
         MCInst2_MC1_r3Inst_XORInst_0_2_n7, MCInst2_MC1_r3Inst_XORInst_0_3_n8,
         MCInst2_MC1_r3Inst_XORInst_0_3_n7, MCInst2_MC2_v1_0_0_,
         MCInst2_MC2_v0_2Inst_0_n3, MCInst2_MC2_v1_2Inst_0_n3,
         MCInst2_MC2_v2_3Inst_0_n6, MCInst2_MC2_v2_3Inst_0_n5,
         MCInst2_MC2_v3_3Inst_0_n3, MCInst2_MC2_v0_2Inst_1_n3,
         MCInst2_MC2_v2_1Inst_1_n3, MCInst2_MC2_v2_2Inst_1_n6,
         MCInst2_MC2_v2_2Inst_1_n5, MCInst2_MC2_v3_3Inst_1_n3,
         MCInst2_MC2_v1_1Inst_2_n3, MCInst2_MC2_v1_2Inst_2_n3,
         MCInst2_MC2_v2_1Inst_2_n3, MCInst2_MC2_v2_2Inst_2_n3,
         MCInst2_MC2_v3_1Inst_2_n3, MCInst2_MC2_v1_2Inst_3_n6,
         MCInst2_MC2_v1_2Inst_3_n5, MCInst2_MC2_v2_2Inst_3_n3,
         MCInst2_MC2_v2_3Inst_3_n3, MCInst2_MC2_r0Inst_XORInst_0_0_n8,
         MCInst2_MC2_r0Inst_XORInst_0_0_n7, MCInst2_MC2_r0Inst_XORInst_0_1_n8,
         MCInst2_MC2_r0Inst_XORInst_0_1_n7, MCInst2_MC2_r0Inst_XORInst_0_2_n8,
         MCInst2_MC2_r0Inst_XORInst_0_2_n7, MCInst2_MC2_r0Inst_XORInst_0_3_n8,
         MCInst2_MC2_r0Inst_XORInst_0_3_n7, MCInst2_MC2_r1Inst_XORInst_0_0_n8,
         MCInst2_MC2_r1Inst_XORInst_0_0_n7, MCInst2_MC2_r1Inst_XORInst_0_1_n8,
         MCInst2_MC2_r1Inst_XORInst_0_1_n7, MCInst2_MC2_r1Inst_XORInst_0_2_n8,
         MCInst2_MC2_r1Inst_XORInst_0_2_n7, MCInst2_MC2_r1Inst_XORInst_0_3_n8,
         MCInst2_MC2_r1Inst_XORInst_0_3_n7, MCInst2_MC2_r2Inst_XORInst_0_0_n8,
         MCInst2_MC2_r2Inst_XORInst_0_0_n7, MCInst2_MC2_r2Inst_XORInst_0_1_n8,
         MCInst2_MC2_r2Inst_XORInst_0_1_n7, MCInst2_MC2_r2Inst_XORInst_0_2_n8,
         MCInst2_MC2_r2Inst_XORInst_0_2_n7, MCInst2_MC2_r2Inst_XORInst_0_3_n8,
         MCInst2_MC2_r2Inst_XORInst_0_3_n7, MCInst2_MC2_r3Inst_XORInst_0_0_n8,
         MCInst2_MC2_r3Inst_XORInst_0_0_n7, MCInst2_MC2_r3Inst_XORInst_0_1_n8,
         MCInst2_MC2_r3Inst_XORInst_0_1_n7, MCInst2_MC2_r3Inst_XORInst_0_2_n8,
         MCInst2_MC2_r3Inst_XORInst_0_2_n7, MCInst2_MC2_r3Inst_XORInst_0_3_n8,
         MCInst2_MC2_r3Inst_XORInst_0_3_n7, MCInst2_MC3_v1_0_0_,
         MCInst2_MC3_v0_2Inst_0_n3, MCInst2_MC3_v1_2Inst_0_n3,
         MCInst2_MC3_v2_3Inst_0_n6, MCInst2_MC3_v2_3Inst_0_n5,
         MCInst2_MC3_v3_3Inst_0_n3, MCInst2_MC3_v0_2Inst_1_n3,
         MCInst2_MC3_v2_1Inst_1_n3, MCInst2_MC3_v2_2Inst_1_n6,
         MCInst2_MC3_v2_2Inst_1_n5, MCInst2_MC3_v3_3Inst_1_n3,
         MCInst2_MC3_v1_1Inst_2_n3, MCInst2_MC3_v1_2Inst_2_n3,
         MCInst2_MC3_v2_1Inst_2_n3, MCInst2_MC3_v2_2Inst_2_n3,
         MCInst2_MC3_v3_1Inst_2_n3, MCInst2_MC3_v1_2Inst_3_n6,
         MCInst2_MC3_v1_2Inst_3_n5, MCInst2_MC3_v2_2Inst_3_n3,
         MCInst2_MC3_v2_3Inst_3_n3, MCInst2_MC3_r0Inst_XORInst_0_0_n8,
         MCInst2_MC3_r0Inst_XORInst_0_0_n7, MCInst2_MC3_r0Inst_XORInst_0_1_n8,
         MCInst2_MC3_r0Inst_XORInst_0_1_n7, MCInst2_MC3_r0Inst_XORInst_0_2_n8,
         MCInst2_MC3_r0Inst_XORInst_0_2_n7, MCInst2_MC3_r0Inst_XORInst_0_3_n8,
         MCInst2_MC3_r0Inst_XORInst_0_3_n7, MCInst2_MC3_r1Inst_XORInst_0_0_n8,
         MCInst2_MC3_r1Inst_XORInst_0_0_n7, MCInst2_MC3_r1Inst_XORInst_0_1_n8,
         MCInst2_MC3_r1Inst_XORInst_0_1_n7, MCInst2_MC3_r1Inst_XORInst_0_2_n8,
         MCInst2_MC3_r1Inst_XORInst_0_2_n7, MCInst2_MC3_r1Inst_XORInst_0_3_n8,
         MCInst2_MC3_r1Inst_XORInst_0_3_n7, MCInst2_MC3_r2Inst_XORInst_0_0_n8,
         MCInst2_MC3_r2Inst_XORInst_0_0_n7, MCInst2_MC3_r2Inst_XORInst_0_1_n8,
         MCInst2_MC3_r2Inst_XORInst_0_1_n7, MCInst2_MC3_r2Inst_XORInst_0_2_n8,
         MCInst2_MC3_r2Inst_XORInst_0_2_n7, MCInst2_MC3_r2Inst_XORInst_0_3_n8,
         MCInst2_MC3_r2Inst_XORInst_0_3_n7, MCInst2_MC3_r3Inst_XORInst_0_0_n8,
         MCInst2_MC3_r3Inst_XORInst_0_0_n7, MCInst2_MC3_r3Inst_XORInst_0_1_n8,
         MCInst2_MC3_r3Inst_XORInst_0_1_n7, MCInst2_MC3_r3Inst_XORInst_0_2_n8,
         MCInst2_MC3_r3Inst_XORInst_0_2_n7, MCInst2_MC3_r3Inst_XORInst_0_3_n8,
         MCInst2_MC3_r3Inst_XORInst_0_3_n7,
         Red_PlaintextInst_LFInst_0_LFInst_0_n3,
         Red_PlaintextInst_LFInst_0_LFInst_1_n3,
         Red_PlaintextInst_LFInst_0_LFInst_2_n3,
         Red_PlaintextInst_LFInst_1_LFInst_0_n3,
         Red_PlaintextInst_LFInst_1_LFInst_1_n3,
         Red_PlaintextInst_LFInst_1_LFInst_2_n3,
         Red_PlaintextInst_LFInst_2_LFInst_0_n3,
         Red_PlaintextInst_LFInst_2_LFInst_1_n3,
         Red_PlaintextInst_LFInst_2_LFInst_2_n3,
         Red_PlaintextInst_LFInst_3_LFInst_0_n3,
         Red_PlaintextInst_LFInst_3_LFInst_1_n3,
         Red_PlaintextInst_LFInst_3_LFInst_2_n3,
         Red_PlaintextInst_LFInst_4_LFInst_0_n3,
         Red_PlaintextInst_LFInst_4_LFInst_1_n3,
         Red_PlaintextInst_LFInst_4_LFInst_2_n3,
         Red_PlaintextInst_LFInst_5_LFInst_0_n3,
         Red_PlaintextInst_LFInst_5_LFInst_1_n3,
         Red_PlaintextInst_LFInst_5_LFInst_2_n3,
         Red_PlaintextInst_LFInst_6_LFInst_0_n3,
         Red_PlaintextInst_LFInst_6_LFInst_1_n3,
         Red_PlaintextInst_LFInst_6_LFInst_2_n3,
         Red_PlaintextInst_LFInst_7_LFInst_0_n3,
         Red_PlaintextInst_LFInst_7_LFInst_1_n3,
         Red_PlaintextInst_LFInst_7_LFInst_2_n3,
         Red_PlaintextInst_LFInst_8_LFInst_0_n3,
         Red_PlaintextInst_LFInst_8_LFInst_1_n3,
         Red_PlaintextInst_LFInst_8_LFInst_2_n3,
         Red_PlaintextInst_LFInst_9_LFInst_0_n3,
         Red_PlaintextInst_LFInst_9_LFInst_1_n3,
         Red_PlaintextInst_LFInst_9_LFInst_2_n3,
         Red_PlaintextInst_LFInst_10_LFInst_0_n3,
         Red_PlaintextInst_LFInst_10_LFInst_1_n3,
         Red_PlaintextInst_LFInst_10_LFInst_2_n3,
         Red_PlaintextInst_LFInst_11_LFInst_0_n3,
         Red_PlaintextInst_LFInst_11_LFInst_1_n3,
         Red_PlaintextInst_LFInst_11_LFInst_2_n3,
         Red_PlaintextInst_LFInst_12_LFInst_0_n3,
         Red_PlaintextInst_LFInst_12_LFInst_1_n3,
         Red_PlaintextInst_LFInst_12_LFInst_2_n3,
         Red_PlaintextInst_LFInst_13_LFInst_0_n3,
         Red_PlaintextInst_LFInst_13_LFInst_1_n3,
         Red_PlaintextInst_LFInst_13_LFInst_2_n3,
         Red_PlaintextInst_LFInst_14_LFInst_0_n3,
         Red_PlaintextInst_LFInst_14_LFInst_1_n3,
         Red_PlaintextInst_LFInst_14_LFInst_2_n3,
         Red_PlaintextInst_LFInst_15_LFInst_0_n3,
         Red_PlaintextInst_LFInst_15_LFInst_1_n3,
         Red_PlaintextInst_LFInst_15_LFInst_2_n3,
         Red_SubCellInst_LFInst_0_LFInst_0_n12,
         Red_SubCellInst_LFInst_0_LFInst_0_n11,
         Red_SubCellInst_LFInst_0_LFInst_0_n10,
         Red_SubCellInst_LFInst_0_LFInst_0_n9,
         Red_SubCellInst_LFInst_0_LFInst_1_n6,
         Red_SubCellInst_LFInst_0_LFInst_1_n5,
         Red_SubCellInst_LFInst_0_LFInst_2_n16,
         Red_SubCellInst_LFInst_0_LFInst_2_n15,
         Red_SubCellInst_LFInst_0_LFInst_2_n14,
         Red_SubCellInst_LFInst_0_LFInst_2_n13,
         Red_SubCellInst_LFInst_0_LFInst_2_n12,
         Red_SubCellInst_LFInst_1_LFInst_0_n12,
         Red_SubCellInst_LFInst_1_LFInst_0_n11,
         Red_SubCellInst_LFInst_1_LFInst_0_n10,
         Red_SubCellInst_LFInst_1_LFInst_0_n9,
         Red_SubCellInst_LFInst_1_LFInst_1_n6,
         Red_SubCellInst_LFInst_1_LFInst_1_n5,
         Red_SubCellInst_LFInst_1_LFInst_2_n16,
         Red_SubCellInst_LFInst_1_LFInst_2_n15,
         Red_SubCellInst_LFInst_1_LFInst_2_n14,
         Red_SubCellInst_LFInst_1_LFInst_2_n13,
         Red_SubCellInst_LFInst_1_LFInst_2_n12,
         Red_SubCellInst_LFInst_2_LFInst_0_n12,
         Red_SubCellInst_LFInst_2_LFInst_0_n11,
         Red_SubCellInst_LFInst_2_LFInst_0_n10,
         Red_SubCellInst_LFInst_2_LFInst_0_n9,
         Red_SubCellInst_LFInst_2_LFInst_1_n6,
         Red_SubCellInst_LFInst_2_LFInst_1_n5,
         Red_SubCellInst_LFInst_2_LFInst_2_n16,
         Red_SubCellInst_LFInst_2_LFInst_2_n15,
         Red_SubCellInst_LFInst_2_LFInst_2_n14,
         Red_SubCellInst_LFInst_2_LFInst_2_n13,
         Red_SubCellInst_LFInst_2_LFInst_2_n12,
         Red_SubCellInst_LFInst_3_LFInst_0_n12,
         Red_SubCellInst_LFInst_3_LFInst_0_n11,
         Red_SubCellInst_LFInst_3_LFInst_0_n10,
         Red_SubCellInst_LFInst_3_LFInst_0_n9,
         Red_SubCellInst_LFInst_3_LFInst_1_n6,
         Red_SubCellInst_LFInst_3_LFInst_1_n5,
         Red_SubCellInst_LFInst_3_LFInst_2_n16,
         Red_SubCellInst_LFInst_3_LFInst_2_n15,
         Red_SubCellInst_LFInst_3_LFInst_2_n14,
         Red_SubCellInst_LFInst_3_LFInst_2_n13,
         Red_SubCellInst_LFInst_3_LFInst_2_n12,
         Red_SubCellInst_LFInst_4_LFInst_0_n12,
         Red_SubCellInst_LFInst_4_LFInst_0_n11,
         Red_SubCellInst_LFInst_4_LFInst_0_n10,
         Red_SubCellInst_LFInst_4_LFInst_0_n9,
         Red_SubCellInst_LFInst_4_LFInst_1_n6,
         Red_SubCellInst_LFInst_4_LFInst_1_n5,
         Red_SubCellInst_LFInst_4_LFInst_2_n16,
         Red_SubCellInst_LFInst_4_LFInst_2_n15,
         Red_SubCellInst_LFInst_4_LFInst_2_n14,
         Red_SubCellInst_LFInst_4_LFInst_2_n13,
         Red_SubCellInst_LFInst_4_LFInst_2_n12,
         Red_SubCellInst_LFInst_5_LFInst_0_n12,
         Red_SubCellInst_LFInst_5_LFInst_0_n11,
         Red_SubCellInst_LFInst_5_LFInst_0_n10,
         Red_SubCellInst_LFInst_5_LFInst_0_n9,
         Red_SubCellInst_LFInst_5_LFInst_1_n6,
         Red_SubCellInst_LFInst_5_LFInst_1_n5,
         Red_SubCellInst_LFInst_5_LFInst_2_n16,
         Red_SubCellInst_LFInst_5_LFInst_2_n15,
         Red_SubCellInst_LFInst_5_LFInst_2_n14,
         Red_SubCellInst_LFInst_5_LFInst_2_n13,
         Red_SubCellInst_LFInst_5_LFInst_2_n12,
         Red_SubCellInst_LFInst_6_LFInst_0_n12,
         Red_SubCellInst_LFInst_6_LFInst_0_n11,
         Red_SubCellInst_LFInst_6_LFInst_0_n10,
         Red_SubCellInst_LFInst_6_LFInst_0_n9,
         Red_SubCellInst_LFInst_6_LFInst_1_n6,
         Red_SubCellInst_LFInst_6_LFInst_1_n5,
         Red_SubCellInst_LFInst_6_LFInst_2_n17,
         Red_SubCellInst_LFInst_6_LFInst_2_n16,
         Red_SubCellInst_LFInst_6_LFInst_2_n15,
         Red_SubCellInst_LFInst_6_LFInst_2_n14,
         Red_SubCellInst_LFInst_6_LFInst_2_n13,
         Red_SubCellInst_LFInst_6_LFInst_2_n12,
         Red_SubCellInst_LFInst_7_LFInst_0_n12,
         Red_SubCellInst_LFInst_7_LFInst_0_n11,
         Red_SubCellInst_LFInst_7_LFInst_0_n10,
         Red_SubCellInst_LFInst_7_LFInst_0_n9,
         Red_SubCellInst_LFInst_7_LFInst_1_n6,
         Red_SubCellInst_LFInst_7_LFInst_1_n5,
         Red_SubCellInst_LFInst_7_LFInst_2_n16,
         Red_SubCellInst_LFInst_7_LFInst_2_n15,
         Red_SubCellInst_LFInst_7_LFInst_2_n14,
         Red_SubCellInst_LFInst_7_LFInst_2_n13,
         Red_SubCellInst_LFInst_7_LFInst_2_n12,
         Red_SubCellInst_LFInst_8_LFInst_0_n12,
         Red_SubCellInst_LFInst_8_LFInst_0_n11,
         Red_SubCellInst_LFInst_8_LFInst_0_n10,
         Red_SubCellInst_LFInst_8_LFInst_0_n9,
         Red_SubCellInst_LFInst_8_LFInst_1_n6,
         Red_SubCellInst_LFInst_8_LFInst_1_n5,
         Red_SubCellInst_LFInst_8_LFInst_2_n13,
         Red_SubCellInst_LFInst_8_LFInst_2_n12,
         Red_SubCellInst_LFInst_8_LFInst_2_n11,
         Red_SubCellInst_LFInst_8_LFInst_2_n10,
         Red_SubCellInst_LFInst_8_LFInst_2_n9,
         Red_SubCellInst_LFInst_9_LFInst_0_n12,
         Red_SubCellInst_LFInst_9_LFInst_0_n11,
         Red_SubCellInst_LFInst_9_LFInst_0_n10,
         Red_SubCellInst_LFInst_9_LFInst_0_n9,
         Red_SubCellInst_LFInst_9_LFInst_1_n6,
         Red_SubCellInst_LFInst_9_LFInst_1_n5,
         Red_SubCellInst_LFInst_9_LFInst_2_n16,
         Red_SubCellInst_LFInst_9_LFInst_2_n15,
         Red_SubCellInst_LFInst_9_LFInst_2_n14,
         Red_SubCellInst_LFInst_9_LFInst_2_n13,
         Red_SubCellInst_LFInst_9_LFInst_2_n12,
         Red_SubCellInst_LFInst_10_LFInst_0_n12,
         Red_SubCellInst_LFInst_10_LFInst_0_n11,
         Red_SubCellInst_LFInst_10_LFInst_0_n10,
         Red_SubCellInst_LFInst_10_LFInst_0_n9,
         Red_SubCellInst_LFInst_10_LFInst_1_n6,
         Red_SubCellInst_LFInst_10_LFInst_1_n5,
         Red_SubCellInst_LFInst_10_LFInst_2_n16,
         Red_SubCellInst_LFInst_10_LFInst_2_n15,
         Red_SubCellInst_LFInst_10_LFInst_2_n14,
         Red_SubCellInst_LFInst_10_LFInst_2_n13,
         Red_SubCellInst_LFInst_10_LFInst_2_n12,
         Red_SubCellInst_LFInst_11_LFInst_0_n12,
         Red_SubCellInst_LFInst_11_LFInst_0_n11,
         Red_SubCellInst_LFInst_11_LFInst_0_n10,
         Red_SubCellInst_LFInst_11_LFInst_0_n9,
         Red_SubCellInst_LFInst_11_LFInst_1_n6,
         Red_SubCellInst_LFInst_11_LFInst_1_n5,
         Red_SubCellInst_LFInst_11_LFInst_2_n16,
         Red_SubCellInst_LFInst_11_LFInst_2_n15,
         Red_SubCellInst_LFInst_11_LFInst_2_n14,
         Red_SubCellInst_LFInst_11_LFInst_2_n13,
         Red_SubCellInst_LFInst_11_LFInst_2_n12,
         Red_SubCellInst_LFInst_12_LFInst_0_n12,
         Red_SubCellInst_LFInst_12_LFInst_0_n11,
         Red_SubCellInst_LFInst_12_LFInst_0_n10,
         Red_SubCellInst_LFInst_12_LFInst_0_n9,
         Red_SubCellInst_LFInst_12_LFInst_1_n6,
         Red_SubCellInst_LFInst_12_LFInst_1_n5,
         Red_SubCellInst_LFInst_12_LFInst_2_n16,
         Red_SubCellInst_LFInst_12_LFInst_2_n15,
         Red_SubCellInst_LFInst_12_LFInst_2_n14,
         Red_SubCellInst_LFInst_12_LFInst_2_n13,
         Red_SubCellInst_LFInst_12_LFInst_2_n12,
         Red_SubCellInst_LFInst_13_LFInst_0_n12,
         Red_SubCellInst_LFInst_13_LFInst_0_n11,
         Red_SubCellInst_LFInst_13_LFInst_0_n10,
         Red_SubCellInst_LFInst_13_LFInst_0_n9,
         Red_SubCellInst_LFInst_13_LFInst_1_n6,
         Red_SubCellInst_LFInst_13_LFInst_1_n5,
         Red_SubCellInst_LFInst_13_LFInst_2_n16,
         Red_SubCellInst_LFInst_13_LFInst_2_n15,
         Red_SubCellInst_LFInst_13_LFInst_2_n14,
         Red_SubCellInst_LFInst_13_LFInst_2_n13,
         Red_SubCellInst_LFInst_13_LFInst_2_n12,
         Red_SubCellInst_LFInst_14_LFInst_0_n12,
         Red_SubCellInst_LFInst_14_LFInst_0_n11,
         Red_SubCellInst_LFInst_14_LFInst_0_n10,
         Red_SubCellInst_LFInst_14_LFInst_0_n9,
         Red_SubCellInst_LFInst_14_LFInst_1_n6,
         Red_SubCellInst_LFInst_14_LFInst_1_n5,
         Red_SubCellInst_LFInst_14_LFInst_2_n16,
         Red_SubCellInst_LFInst_14_LFInst_2_n15,
         Red_SubCellInst_LFInst_14_LFInst_2_n14,
         Red_SubCellInst_LFInst_14_LFInst_2_n13,
         Red_SubCellInst_LFInst_14_LFInst_2_n12,
         Red_SubCellInst_LFInst_15_LFInst_0_n12,
         Red_SubCellInst_LFInst_15_LFInst_0_n11,
         Red_SubCellInst_LFInst_15_LFInst_0_n10,
         Red_SubCellInst_LFInst_15_LFInst_0_n9,
         Red_SubCellInst_LFInst_15_LFInst_1_n6,
         Red_SubCellInst_LFInst_15_LFInst_1_n5,
         Red_SubCellInst_LFInst_15_LFInst_2_n16,
         Red_SubCellInst_LFInst_15_LFInst_2_n15,
         Red_SubCellInst_LFInst_15_LFInst_2_n14,
         Red_SubCellInst_LFInst_15_LFInst_2_n13,
         Red_SubCellInst_LFInst_15_LFInst_2_n12, Red_MCInst_MC0_v1_0Inst_0_n3,
         Red_MCInst_MC0_v2_2Inst_0_n3, Red_MCInst_MC0_v2_3Inst_0_n3,
         Red_MCInst_MC0_v3_2Inst_0_n6, Red_MCInst_MC0_v3_2Inst_0_n5,
         Red_MCInst_MC0_v0_1Inst_1_n3, Red_MCInst_MC0_v1_0Inst_1_n3,
         Red_MCInst_MC0_v1_1Inst_1_n6, Red_MCInst_MC0_v1_1Inst_1_n5,
         Red_MCInst_MC0_v3_1Inst_1_n6, Red_MCInst_MC0_v3_1Inst_1_n5,
         Red_MCInst_MC0_v0_0Inst_2_n3, Red_MCInst_MC0_v0_3Inst_2_n6,
         Red_MCInst_MC0_v0_3Inst_2_n5, Red_MCInst_MC0_v1_0Inst_2_n3,
         Red_MCInst_MC0_v1_2Inst_2_n3, Red_MCInst_MC0_v1_3Inst_2_n6,
         Red_MCInst_MC0_v1_3Inst_2_n5, Red_MCInst_MC0_v2_0Inst_2_n6,
         Red_MCInst_MC0_v2_0Inst_2_n5, Red_MCInst_MC0_v3_0Inst_2_n6,
         Red_MCInst_MC0_v3_0Inst_2_n5, Red_MCInst_MC0_v3_2Inst_2_n3,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC0_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC0_r3Inst_XORInst_0_2_n7, Red_MCInst_MC1_v1_0Inst_0_n3,
         Red_MCInst_MC1_v2_2Inst_0_n3, Red_MCInst_MC1_v2_3Inst_0_n3,
         Red_MCInst_MC1_v3_2Inst_0_n6, Red_MCInst_MC1_v3_2Inst_0_n5,
         Red_MCInst_MC1_v0_1Inst_1_n3, Red_MCInst_MC1_v1_0Inst_1_n3,
         Red_MCInst_MC1_v1_1Inst_1_n6, Red_MCInst_MC1_v1_1Inst_1_n5,
         Red_MCInst_MC1_v3_1Inst_1_n6, Red_MCInst_MC1_v3_1Inst_1_n5,
         Red_MCInst_MC1_v0_0Inst_2_n3, Red_MCInst_MC1_v0_3Inst_2_n6,
         Red_MCInst_MC1_v0_3Inst_2_n5, Red_MCInst_MC1_v1_0Inst_2_n3,
         Red_MCInst_MC1_v1_2Inst_2_n3, Red_MCInst_MC1_v1_3Inst_2_n6,
         Red_MCInst_MC1_v1_3Inst_2_n5, Red_MCInst_MC1_v2_0Inst_2_n6,
         Red_MCInst_MC1_v2_0Inst_2_n5, Red_MCInst_MC1_v3_0Inst_2_n6,
         Red_MCInst_MC1_v3_0Inst_2_n5, Red_MCInst_MC1_v3_2Inst_2_n3,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC1_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC1_r3Inst_XORInst_0_2_n7, Red_MCInst_MC2_v1_0Inst_0_n3,
         Red_MCInst_MC2_v2_2Inst_0_n3, Red_MCInst_MC2_v2_3Inst_0_n3,
         Red_MCInst_MC2_v3_2Inst_0_n6, Red_MCInst_MC2_v3_2Inst_0_n5,
         Red_MCInst_MC2_v0_1Inst_1_n3, Red_MCInst_MC2_v1_0Inst_1_n3,
         Red_MCInst_MC2_v1_1Inst_1_n6, Red_MCInst_MC2_v1_1Inst_1_n5,
         Red_MCInst_MC2_v3_1Inst_1_n6, Red_MCInst_MC2_v3_1Inst_1_n5,
         Red_MCInst_MC2_v0_0Inst_2_n3, Red_MCInst_MC2_v0_3Inst_2_n6,
         Red_MCInst_MC2_v0_3Inst_2_n5, Red_MCInst_MC2_v1_0Inst_2_n3,
         Red_MCInst_MC2_v1_2Inst_2_n3, Red_MCInst_MC2_v1_3Inst_2_n6,
         Red_MCInst_MC2_v1_3Inst_2_n5, Red_MCInst_MC2_v2_0Inst_2_n6,
         Red_MCInst_MC2_v2_0Inst_2_n5, Red_MCInst_MC2_v3_0Inst_2_n6,
         Red_MCInst_MC2_v3_0Inst_2_n5, Red_MCInst_MC2_v3_2Inst_2_n3,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC2_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC2_r3Inst_XORInst_0_2_n7, Red_MCInst_MC3_v1_0Inst_0_n3,
         Red_MCInst_MC3_v2_2Inst_0_n3, Red_MCInst_MC3_v2_3Inst_0_n3,
         Red_MCInst_MC3_v3_2Inst_0_n6, Red_MCInst_MC3_v3_2Inst_0_n5,
         Red_MCInst_MC3_v0_1Inst_1_n3, Red_MCInst_MC3_v1_0Inst_1_n3,
         Red_MCInst_MC3_v1_1Inst_1_n6, Red_MCInst_MC3_v1_1Inst_1_n5,
         Red_MCInst_MC3_v3_1Inst_1_n6, Red_MCInst_MC3_v3_1Inst_1_n5,
         Red_MCInst_MC3_v0_0Inst_2_n3, Red_MCInst_MC3_v0_3Inst_2_n6,
         Red_MCInst_MC3_v0_3Inst_2_n5, Red_MCInst_MC3_v1_0Inst_2_n3,
         Red_MCInst_MC3_v1_2Inst_2_n3, Red_MCInst_MC3_v1_3Inst_2_n6,
         Red_MCInst_MC3_v1_3Inst_2_n5, Red_MCInst_MC3_v2_0Inst_2_n6,
         Red_MCInst_MC3_v2_0Inst_2_n5, Red_MCInst_MC3_v3_0Inst_2_n6,
         Red_MCInst_MC3_v3_0Inst_2_n5, Red_MCInst_MC3_v3_2Inst_2_n3,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r0Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r0Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r0Inst_XORInst_0_2_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r1Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r1Inst_XORInst_0_2_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r2Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r2Inst_XORInst_0_2_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_1_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_1_n7,
         Red_MCInst_MC3_r3Inst_XORInst_0_2_n8,
         Red_MCInst_MC3_r3Inst_XORInst_0_2_n7,
         Red_SubCellInst2_LFInst_0_LFInst_0_n12,
         Red_SubCellInst2_LFInst_0_LFInst_0_n11,
         Red_SubCellInst2_LFInst_0_LFInst_0_n10,
         Red_SubCellInst2_LFInst_0_LFInst_0_n9,
         Red_SubCellInst2_LFInst_0_LFInst_1_n6,
         Red_SubCellInst2_LFInst_0_LFInst_1_n5,
         Red_SubCellInst2_LFInst_0_LFInst_2_n17,
         Red_SubCellInst2_LFInst_0_LFInst_2_n16,
         Red_SubCellInst2_LFInst_0_LFInst_2_n15,
         Red_SubCellInst2_LFInst_0_LFInst_2_n14,
         Red_SubCellInst2_LFInst_0_LFInst_2_n13,
         Red_SubCellInst2_LFInst_0_LFInst_2_n12,
         Red_SubCellInst2_LFInst_1_LFInst_0_n12,
         Red_SubCellInst2_LFInst_1_LFInst_0_n11,
         Red_SubCellInst2_LFInst_1_LFInst_0_n10,
         Red_SubCellInst2_LFInst_1_LFInst_0_n9,
         Red_SubCellInst2_LFInst_1_LFInst_1_n6,
         Red_SubCellInst2_LFInst_1_LFInst_1_n5,
         Red_SubCellInst2_LFInst_1_LFInst_2_n14,
         Red_SubCellInst2_LFInst_1_LFInst_2_n13,
         Red_SubCellInst2_LFInst_1_LFInst_2_n12,
         Red_SubCellInst2_LFInst_1_LFInst_2_n11,
         Red_SubCellInst2_LFInst_1_LFInst_2_n10,
         Red_SubCellInst2_LFInst_1_LFInst_2_n9,
         Red_SubCellInst2_LFInst_2_LFInst_0_n12,
         Red_SubCellInst2_LFInst_2_LFInst_0_n11,
         Red_SubCellInst2_LFInst_2_LFInst_0_n10,
         Red_SubCellInst2_LFInst_2_LFInst_0_n9,
         Red_SubCellInst2_LFInst_2_LFInst_1_n6,
         Red_SubCellInst2_LFInst_2_LFInst_1_n5,
         Red_SubCellInst2_LFInst_2_LFInst_2_n17,
         Red_SubCellInst2_LFInst_2_LFInst_2_n16,
         Red_SubCellInst2_LFInst_2_LFInst_2_n15,
         Red_SubCellInst2_LFInst_2_LFInst_2_n14,
         Red_SubCellInst2_LFInst_2_LFInst_2_n13,
         Red_SubCellInst2_LFInst_2_LFInst_2_n12,
         Red_SubCellInst2_LFInst_3_LFInst_0_n12,
         Red_SubCellInst2_LFInst_3_LFInst_0_n11,
         Red_SubCellInst2_LFInst_3_LFInst_0_n10,
         Red_SubCellInst2_LFInst_3_LFInst_0_n9,
         Red_SubCellInst2_LFInst_3_LFInst_1_n6,
         Red_SubCellInst2_LFInst_3_LFInst_1_n5,
         Red_SubCellInst2_LFInst_3_LFInst_2_n17,
         Red_SubCellInst2_LFInst_3_LFInst_2_n16,
         Red_SubCellInst2_LFInst_3_LFInst_2_n15,
         Red_SubCellInst2_LFInst_3_LFInst_2_n14,
         Red_SubCellInst2_LFInst_3_LFInst_2_n13,
         Red_SubCellInst2_LFInst_3_LFInst_2_n12,
         Red_SubCellInst2_LFInst_4_LFInst_0_n12,
         Red_SubCellInst2_LFInst_4_LFInst_0_n11,
         Red_SubCellInst2_LFInst_4_LFInst_0_n10,
         Red_SubCellInst2_LFInst_4_LFInst_0_n9,
         Red_SubCellInst2_LFInst_4_LFInst_1_n6,
         Red_SubCellInst2_LFInst_4_LFInst_1_n5,
         Red_SubCellInst2_LFInst_4_LFInst_2_n16,
         Red_SubCellInst2_LFInst_4_LFInst_2_n15,
         Red_SubCellInst2_LFInst_4_LFInst_2_n14,
         Red_SubCellInst2_LFInst_4_LFInst_2_n13,
         Red_SubCellInst2_LFInst_4_LFInst_2_n12,
         Red_SubCellInst2_LFInst_5_LFInst_0_n12,
         Red_SubCellInst2_LFInst_5_LFInst_0_n11,
         Red_SubCellInst2_LFInst_5_LFInst_0_n10,
         Red_SubCellInst2_LFInst_5_LFInst_0_n9,
         Red_SubCellInst2_LFInst_5_LFInst_1_n6,
         Red_SubCellInst2_LFInst_5_LFInst_1_n5,
         Red_SubCellInst2_LFInst_5_LFInst_2_n17,
         Red_SubCellInst2_LFInst_5_LFInst_2_n16,
         Red_SubCellInst2_LFInst_5_LFInst_2_n15,
         Red_SubCellInst2_LFInst_5_LFInst_2_n14,
         Red_SubCellInst2_LFInst_5_LFInst_2_n13,
         Red_SubCellInst2_LFInst_5_LFInst_2_n12,
         Red_SubCellInst2_LFInst_6_LFInst_0_n12,
         Red_SubCellInst2_LFInst_6_LFInst_0_n11,
         Red_SubCellInst2_LFInst_6_LFInst_0_n10,
         Red_SubCellInst2_LFInst_6_LFInst_0_n9,
         Red_SubCellInst2_LFInst_6_LFInst_1_n6,
         Red_SubCellInst2_LFInst_6_LFInst_1_n5,
         Red_SubCellInst2_LFInst_6_LFInst_2_n17,
         Red_SubCellInst2_LFInst_6_LFInst_2_n16,
         Red_SubCellInst2_LFInst_6_LFInst_2_n15,
         Red_SubCellInst2_LFInst_6_LFInst_2_n14,
         Red_SubCellInst2_LFInst_6_LFInst_2_n13,
         Red_SubCellInst2_LFInst_6_LFInst_2_n12,
         Red_SubCellInst2_LFInst_7_LFInst_0_n12,
         Red_SubCellInst2_LFInst_7_LFInst_0_n11,
         Red_SubCellInst2_LFInst_7_LFInst_0_n10,
         Red_SubCellInst2_LFInst_7_LFInst_0_n9,
         Red_SubCellInst2_LFInst_7_LFInst_1_n6,
         Red_SubCellInst2_LFInst_7_LFInst_1_n5,
         Red_SubCellInst2_LFInst_7_LFInst_2_n17,
         Red_SubCellInst2_LFInst_7_LFInst_2_n16,
         Red_SubCellInst2_LFInst_7_LFInst_2_n15,
         Red_SubCellInst2_LFInst_7_LFInst_2_n14,
         Red_SubCellInst2_LFInst_7_LFInst_2_n13,
         Red_SubCellInst2_LFInst_7_LFInst_2_n12,
         Red_SubCellInst2_LFInst_8_LFInst_0_n12,
         Red_SubCellInst2_LFInst_8_LFInst_0_n11,
         Red_SubCellInst2_LFInst_8_LFInst_0_n10,
         Red_SubCellInst2_LFInst_8_LFInst_0_n9,
         Red_SubCellInst2_LFInst_8_LFInst_1_n6,
         Red_SubCellInst2_LFInst_8_LFInst_1_n5,
         Red_SubCellInst2_LFInst_8_LFInst_2_n14,
         Red_SubCellInst2_LFInst_8_LFInst_2_n13,
         Red_SubCellInst2_LFInst_8_LFInst_2_n12,
         Red_SubCellInst2_LFInst_8_LFInst_2_n11,
         Red_SubCellInst2_LFInst_8_LFInst_2_n10,
         Red_SubCellInst2_LFInst_8_LFInst_2_n9,
         Red_SubCellInst2_LFInst_9_LFInst_0_n12,
         Red_SubCellInst2_LFInst_9_LFInst_0_n11,
         Red_SubCellInst2_LFInst_9_LFInst_0_n10,
         Red_SubCellInst2_LFInst_9_LFInst_0_n9,
         Red_SubCellInst2_LFInst_9_LFInst_1_n6,
         Red_SubCellInst2_LFInst_9_LFInst_1_n5,
         Red_SubCellInst2_LFInst_9_LFInst_2_n16,
         Red_SubCellInst2_LFInst_9_LFInst_2_n15,
         Red_SubCellInst2_LFInst_9_LFInst_2_n14,
         Red_SubCellInst2_LFInst_9_LFInst_2_n13,
         Red_SubCellInst2_LFInst_9_LFInst_2_n12,
         Red_SubCellInst2_LFInst_10_LFInst_0_n12,
         Red_SubCellInst2_LFInst_10_LFInst_0_n11,
         Red_SubCellInst2_LFInst_10_LFInst_0_n10,
         Red_SubCellInst2_LFInst_10_LFInst_0_n9,
         Red_SubCellInst2_LFInst_10_LFInst_1_n6,
         Red_SubCellInst2_LFInst_10_LFInst_1_n5,
         Red_SubCellInst2_LFInst_10_LFInst_2_n17,
         Red_SubCellInst2_LFInst_10_LFInst_2_n16,
         Red_SubCellInst2_LFInst_10_LFInst_2_n15,
         Red_SubCellInst2_LFInst_10_LFInst_2_n14,
         Red_SubCellInst2_LFInst_10_LFInst_2_n13,
         Red_SubCellInst2_LFInst_10_LFInst_2_n12,
         Red_SubCellInst2_LFInst_11_LFInst_0_n12,
         Red_SubCellInst2_LFInst_11_LFInst_0_n11,
         Red_SubCellInst2_LFInst_11_LFInst_0_n10,
         Red_SubCellInst2_LFInst_11_LFInst_0_n9,
         Red_SubCellInst2_LFInst_11_LFInst_1_n6,
         Red_SubCellInst2_LFInst_11_LFInst_1_n5,
         Red_SubCellInst2_LFInst_11_LFInst_2_n17,
         Red_SubCellInst2_LFInst_11_LFInst_2_n16,
         Red_SubCellInst2_LFInst_11_LFInst_2_n15,
         Red_SubCellInst2_LFInst_11_LFInst_2_n14,
         Red_SubCellInst2_LFInst_11_LFInst_2_n13,
         Red_SubCellInst2_LFInst_11_LFInst_2_n12,
         Red_SubCellInst2_LFInst_12_LFInst_0_n12,
         Red_SubCellInst2_LFInst_12_LFInst_0_n11,
         Red_SubCellInst2_LFInst_12_LFInst_0_n10,
         Red_SubCellInst2_LFInst_12_LFInst_0_n9,
         Red_SubCellInst2_LFInst_12_LFInst_1_n6,
         Red_SubCellInst2_LFInst_12_LFInst_1_n5,
         Red_SubCellInst2_LFInst_12_LFInst_2_n16,
         Red_SubCellInst2_LFInst_12_LFInst_2_n15,
         Red_SubCellInst2_LFInst_12_LFInst_2_n14,
         Red_SubCellInst2_LFInst_12_LFInst_2_n13,
         Red_SubCellInst2_LFInst_12_LFInst_2_n12,
         Red_SubCellInst2_LFInst_13_LFInst_0_n12,
         Red_SubCellInst2_LFInst_13_LFInst_0_n11,
         Red_SubCellInst2_LFInst_13_LFInst_0_n10,
         Red_SubCellInst2_LFInst_13_LFInst_0_n9,
         Red_SubCellInst2_LFInst_13_LFInst_1_n6,
         Red_SubCellInst2_LFInst_13_LFInst_1_n5,
         Red_SubCellInst2_LFInst_13_LFInst_2_n17,
         Red_SubCellInst2_LFInst_13_LFInst_2_n16,
         Red_SubCellInst2_LFInst_13_LFInst_2_n15,
         Red_SubCellInst2_LFInst_13_LFInst_2_n14,
         Red_SubCellInst2_LFInst_13_LFInst_2_n13,
         Red_SubCellInst2_LFInst_13_LFInst_2_n12,
         Red_SubCellInst2_LFInst_14_LFInst_0_n12,
         Red_SubCellInst2_LFInst_14_LFInst_0_n11,
         Red_SubCellInst2_LFInst_14_LFInst_0_n10,
         Red_SubCellInst2_LFInst_14_LFInst_0_n9,
         Red_SubCellInst2_LFInst_14_LFInst_1_n6,
         Red_SubCellInst2_LFInst_14_LFInst_1_n5,
         Red_SubCellInst2_LFInst_14_LFInst_2_n16,
         Red_SubCellInst2_LFInst_14_LFInst_2_n15,
         Red_SubCellInst2_LFInst_14_LFInst_2_n14,
         Red_SubCellInst2_LFInst_14_LFInst_2_n13,
         Red_SubCellInst2_LFInst_14_LFInst_2_n12,
         Red_SubCellInst2_LFInst_15_LFInst_0_n12,
         Red_SubCellInst2_LFInst_15_LFInst_0_n11,
         Red_SubCellInst2_LFInst_15_LFInst_0_n10,
         Red_SubCellInst2_LFInst_15_LFInst_0_n9,
         Red_SubCellInst2_LFInst_15_LFInst_1_n6,
         Red_SubCellInst2_LFInst_15_LFInst_1_n5,
         Red_SubCellInst2_LFInst_15_LFInst_2_n17,
         Red_SubCellInst2_LFInst_15_LFInst_2_n16,
         Red_SubCellInst2_LFInst_15_LFInst_2_n15,
         Red_SubCellInst2_LFInst_15_LFInst_2_n14,
         Red_SubCellInst2_LFInst_15_LFInst_2_n13,
         Red_SubCellInst2_LFInst_15_LFInst_2_n12,
         Red_MCInst2_MC0_v1_0Inst_0_n3, Red_MCInst2_MC0_v2_2Inst_0_n3,
         Red_MCInst2_MC0_v2_3Inst_0_n3, Red_MCInst2_MC0_v3_2Inst_0_n6,
         Red_MCInst2_MC0_v3_2Inst_0_n5, Red_MCInst2_MC0_v0_1Inst_1_n3,
         Red_MCInst2_MC0_v1_0Inst_1_n3, Red_MCInst2_MC0_v1_1Inst_1_n6,
         Red_MCInst2_MC0_v1_1Inst_1_n5, Red_MCInst2_MC0_v3_1Inst_1_n6,
         Red_MCInst2_MC0_v3_1Inst_1_n5, Red_MCInst2_MC0_v0_0Inst_2_n3,
         Red_MCInst2_MC0_v0_3Inst_2_n6, Red_MCInst2_MC0_v0_3Inst_2_n5,
         Red_MCInst2_MC0_v1_0Inst_2_n3, Red_MCInst2_MC0_v1_2Inst_2_n3,
         Red_MCInst2_MC0_v1_3Inst_2_n6, Red_MCInst2_MC0_v1_3Inst_2_n5,
         Red_MCInst2_MC0_v2_0Inst_2_n6, Red_MCInst2_MC0_v2_0Inst_2_n5,
         Red_MCInst2_MC0_v3_0Inst_2_n6, Red_MCInst2_MC0_v3_0Inst_2_n5,
         Red_MCInst2_MC0_v3_2Inst_2_n3, Red_MCInst2_MC0_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r0Inst_XORInst_0_1_n8,
         Red_MCInst2_MC0_r0Inst_XORInst_0_1_n7,
         Red_MCInst2_MC0_r0Inst_XORInst_0_2_n8,
         Red_MCInst2_MC0_r0Inst_XORInst_0_2_n7,
         Red_MCInst2_MC0_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r1Inst_XORInst_0_1_n8,
         Red_MCInst2_MC0_r1Inst_XORInst_0_1_n7,
         Red_MCInst2_MC0_r1Inst_XORInst_0_2_n8,
         Red_MCInst2_MC0_r1Inst_XORInst_0_2_n7,
         Red_MCInst2_MC0_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r2Inst_XORInst_0_1_n8,
         Red_MCInst2_MC0_r2Inst_XORInst_0_1_n7,
         Red_MCInst2_MC0_r2Inst_XORInst_0_2_n8,
         Red_MCInst2_MC0_r2Inst_XORInst_0_2_n7,
         Red_MCInst2_MC0_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC0_r3Inst_XORInst_0_0_n7,
         Red_MCInst2_MC0_r3Inst_XORInst_0_1_n8,
         Red_MCInst2_MC0_r3Inst_XORInst_0_1_n7,
         Red_MCInst2_MC0_r3Inst_XORInst_0_2_n8,
         Red_MCInst2_MC0_r3Inst_XORInst_0_2_n7, Red_MCInst2_MC1_v1_0Inst_0_n3,
         Red_MCInst2_MC1_v2_2Inst_0_n3, Red_MCInst2_MC1_v2_3Inst_0_n3,
         Red_MCInst2_MC1_v3_2Inst_0_n6, Red_MCInst2_MC1_v3_2Inst_0_n5,
         Red_MCInst2_MC1_v0_1Inst_1_n3, Red_MCInst2_MC1_v1_0Inst_1_n3,
         Red_MCInst2_MC1_v1_1Inst_1_n6, Red_MCInst2_MC1_v1_1Inst_1_n5,
         Red_MCInst2_MC1_v3_1Inst_1_n6, Red_MCInst2_MC1_v3_1Inst_1_n5,
         Red_MCInst2_MC1_v0_0Inst_2_n3, Red_MCInst2_MC1_v0_3Inst_2_n6,
         Red_MCInst2_MC1_v0_3Inst_2_n5, Red_MCInst2_MC1_v1_0Inst_2_n3,
         Red_MCInst2_MC1_v1_2Inst_2_n3, Red_MCInst2_MC1_v1_3Inst_2_n6,
         Red_MCInst2_MC1_v1_3Inst_2_n5, Red_MCInst2_MC1_v2_0Inst_2_n6,
         Red_MCInst2_MC1_v2_0Inst_2_n5, Red_MCInst2_MC1_v3_0Inst_2_n6,
         Red_MCInst2_MC1_v3_0Inst_2_n5, Red_MCInst2_MC1_v3_2Inst_2_n3,
         Red_MCInst2_MC1_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r0Inst_XORInst_0_1_n8,
         Red_MCInst2_MC1_r0Inst_XORInst_0_1_n7,
         Red_MCInst2_MC1_r0Inst_XORInst_0_2_n8,
         Red_MCInst2_MC1_r0Inst_XORInst_0_2_n7,
         Red_MCInst2_MC1_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r1Inst_XORInst_0_1_n8,
         Red_MCInst2_MC1_r1Inst_XORInst_0_1_n7,
         Red_MCInst2_MC1_r1Inst_XORInst_0_2_n8,
         Red_MCInst2_MC1_r1Inst_XORInst_0_2_n7,
         Red_MCInst2_MC1_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r2Inst_XORInst_0_1_n8,
         Red_MCInst2_MC1_r2Inst_XORInst_0_1_n7,
         Red_MCInst2_MC1_r2Inst_XORInst_0_2_n8,
         Red_MCInst2_MC1_r2Inst_XORInst_0_2_n7,
         Red_MCInst2_MC1_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC1_r3Inst_XORInst_0_0_n7,
         Red_MCInst2_MC1_r3Inst_XORInst_0_1_n8,
         Red_MCInst2_MC1_r3Inst_XORInst_0_1_n7,
         Red_MCInst2_MC1_r3Inst_XORInst_0_2_n8,
         Red_MCInst2_MC1_r3Inst_XORInst_0_2_n7, Red_MCInst2_MC2_v1_0Inst_0_n3,
         Red_MCInst2_MC2_v2_2Inst_0_n3, Red_MCInst2_MC2_v2_3Inst_0_n3,
         Red_MCInst2_MC2_v3_2Inst_0_n6, Red_MCInst2_MC2_v3_2Inst_0_n5,
         Red_MCInst2_MC2_v0_1Inst_1_n3, Red_MCInst2_MC2_v1_0Inst_1_n3,
         Red_MCInst2_MC2_v1_1Inst_1_n6, Red_MCInst2_MC2_v1_1Inst_1_n5,
         Red_MCInst2_MC2_v3_1Inst_1_n6, Red_MCInst2_MC2_v3_1Inst_1_n5,
         Red_MCInst2_MC2_v0_0Inst_2_n3, Red_MCInst2_MC2_v0_3Inst_2_n6,
         Red_MCInst2_MC2_v0_3Inst_2_n5, Red_MCInst2_MC2_v1_0Inst_2_n3,
         Red_MCInst2_MC2_v1_2Inst_2_n3, Red_MCInst2_MC2_v1_3Inst_2_n6,
         Red_MCInst2_MC2_v1_3Inst_2_n5, Red_MCInst2_MC2_v2_0Inst_2_n6,
         Red_MCInst2_MC2_v2_0Inst_2_n5, Red_MCInst2_MC2_v3_0Inst_2_n6,
         Red_MCInst2_MC2_v3_0Inst_2_n5, Red_MCInst2_MC2_v3_2Inst_2_n3,
         Red_MCInst2_MC2_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r0Inst_XORInst_0_1_n8,
         Red_MCInst2_MC2_r0Inst_XORInst_0_1_n7,
         Red_MCInst2_MC2_r0Inst_XORInst_0_2_n8,
         Red_MCInst2_MC2_r0Inst_XORInst_0_2_n7,
         Red_MCInst2_MC2_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r1Inst_XORInst_0_1_n8,
         Red_MCInst2_MC2_r1Inst_XORInst_0_1_n7,
         Red_MCInst2_MC2_r1Inst_XORInst_0_2_n8,
         Red_MCInst2_MC2_r1Inst_XORInst_0_2_n7,
         Red_MCInst2_MC2_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r2Inst_XORInst_0_1_n8,
         Red_MCInst2_MC2_r2Inst_XORInst_0_1_n7,
         Red_MCInst2_MC2_r2Inst_XORInst_0_2_n8,
         Red_MCInst2_MC2_r2Inst_XORInst_0_2_n7,
         Red_MCInst2_MC2_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC2_r3Inst_XORInst_0_0_n7,
         Red_MCInst2_MC2_r3Inst_XORInst_0_1_n8,
         Red_MCInst2_MC2_r3Inst_XORInst_0_1_n7,
         Red_MCInst2_MC2_r3Inst_XORInst_0_2_n8,
         Red_MCInst2_MC2_r3Inst_XORInst_0_2_n7, Red_MCInst2_MC3_v1_0Inst_0_n3,
         Red_MCInst2_MC3_v2_2Inst_0_n3, Red_MCInst2_MC3_v2_3Inst_0_n3,
         Red_MCInst2_MC3_v3_2Inst_0_n6, Red_MCInst2_MC3_v3_2Inst_0_n5,
         Red_MCInst2_MC3_v0_1Inst_1_n3, Red_MCInst2_MC3_v1_0Inst_1_n3,
         Red_MCInst2_MC3_v1_1Inst_1_n6, Red_MCInst2_MC3_v1_1Inst_1_n5,
         Red_MCInst2_MC3_v3_1Inst_1_n6, Red_MCInst2_MC3_v3_1Inst_1_n5,
         Red_MCInst2_MC3_v0_0Inst_2_n3, Red_MCInst2_MC3_v0_3Inst_2_n6,
         Red_MCInst2_MC3_v0_3Inst_2_n5, Red_MCInst2_MC3_v1_0Inst_2_n3,
         Red_MCInst2_MC3_v1_2Inst_2_n3, Red_MCInst2_MC3_v1_3Inst_2_n6,
         Red_MCInst2_MC3_v1_3Inst_2_n5, Red_MCInst2_MC3_v2_0Inst_2_n6,
         Red_MCInst2_MC3_v2_0Inst_2_n5, Red_MCInst2_MC3_v3_0Inst_2_n6,
         Red_MCInst2_MC3_v3_0Inst_2_n5, Red_MCInst2_MC3_v3_2Inst_2_n3,
         Red_MCInst2_MC3_r0Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r0Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r0Inst_XORInst_0_1_n8,
         Red_MCInst2_MC3_r0Inst_XORInst_0_1_n7,
         Red_MCInst2_MC3_r0Inst_XORInst_0_2_n8,
         Red_MCInst2_MC3_r0Inst_XORInst_0_2_n7,
         Red_MCInst2_MC3_r1Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r1Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r1Inst_XORInst_0_1_n8,
         Red_MCInst2_MC3_r1Inst_XORInst_0_1_n7,
         Red_MCInst2_MC3_r1Inst_XORInst_0_2_n8,
         Red_MCInst2_MC3_r1Inst_XORInst_0_2_n7,
         Red_MCInst2_MC3_r2Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r2Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r2Inst_XORInst_0_1_n8,
         Red_MCInst2_MC3_r2Inst_XORInst_0_1_n7,
         Red_MCInst2_MC3_r2Inst_XORInst_0_2_n8,
         Red_MCInst2_MC3_r2Inst_XORInst_0_2_n7,
         Red_MCInst2_MC3_r3Inst_XORInst_0_0_n8,
         Red_MCInst2_MC3_r3Inst_XORInst_0_0_n7,
         Red_MCInst2_MC3_r3Inst_XORInst_0_1_n8,
         Red_MCInst2_MC3_r3Inst_XORInst_0_1_n7,
         Red_MCInst2_MC3_r3Inst_XORInst_0_2_n8,
         Red_MCInst2_MC3_r3Inst_XORInst_0_2_n7,
         Red_KeyInst_LFInst_0_LFInst_0_n3, Red_KeyInst_LFInst_0_LFInst_1_n3,
         Red_KeyInst_LFInst_0_LFInst_2_n3, Red_KeyInst_LFInst_1_LFInst_0_n3,
         Red_KeyInst_LFInst_1_LFInst_1_n3, Red_KeyInst_LFInst_1_LFInst_2_n3,
         Red_KeyInst_LFInst_2_LFInst_0_n3, Red_KeyInst_LFInst_2_LFInst_1_n3,
         Red_KeyInst_LFInst_2_LFInst_2_n3, Red_KeyInst_LFInst_3_LFInst_0_n3,
         Red_KeyInst_LFInst_3_LFInst_1_n3, Red_KeyInst_LFInst_3_LFInst_2_n3,
         Red_KeyInst_LFInst_4_LFInst_0_n3, Red_KeyInst_LFInst_4_LFInst_1_n3,
         Red_KeyInst_LFInst_4_LFInst_2_n3, Red_KeyInst_LFInst_5_LFInst_0_n3,
         Red_KeyInst_LFInst_5_LFInst_1_n3, Red_KeyInst_LFInst_5_LFInst_2_n3,
         Red_KeyInst_LFInst_6_LFInst_0_n3, Red_KeyInst_LFInst_6_LFInst_1_n3,
         Red_KeyInst_LFInst_6_LFInst_2_n3, Red_KeyInst_LFInst_7_LFInst_0_n3,
         Red_KeyInst_LFInst_7_LFInst_1_n3, Red_KeyInst_LFInst_7_LFInst_2_n3,
         Red_KeyInst_LFInst_8_LFInst_0_n3, Red_KeyInst_LFInst_8_LFInst_1_n3,
         Red_KeyInst_LFInst_8_LFInst_2_n3, Red_KeyInst_LFInst_9_LFInst_0_n3,
         Red_KeyInst_LFInst_9_LFInst_1_n3, Red_KeyInst_LFInst_9_LFInst_2_n3,
         Red_KeyInst_LFInst_10_LFInst_0_n3, Red_KeyInst_LFInst_10_LFInst_1_n3,
         Red_KeyInst_LFInst_10_LFInst_2_n3, Red_KeyInst_LFInst_11_LFInst_0_n3,
         Red_KeyInst_LFInst_11_LFInst_1_n3, Red_KeyInst_LFInst_11_LFInst_2_n3,
         Red_KeyInst_LFInst_12_LFInst_0_n3, Red_KeyInst_LFInst_12_LFInst_1_n3,
         Red_KeyInst_LFInst_12_LFInst_2_n3, Red_KeyInst_LFInst_13_LFInst_0_n3,
         Red_KeyInst_LFInst_13_LFInst_1_n3, Red_KeyInst_LFInst_13_LFInst_2_n3,
         Red_KeyInst_LFInst_14_LFInst_0_n3, Red_KeyInst_LFInst_14_LFInst_1_n3,
         Red_KeyInst_LFInst_14_LFInst_2_n3, Red_KeyInst_LFInst_15_LFInst_0_n3,
         Red_KeyInst_LFInst_15_LFInst_1_n3, Red_KeyInst_LFInst_15_LFInst_2_n3,
         Red_ToCheckInst_LFInst_0_LFInst_0_n3,
         Red_ToCheckInst_LFInst_0_LFInst_1_n3,
         Red_ToCheckInst_LFInst_0_LFInst_2_n3,
         Red_ToCheckInst_LFInst_1_LFInst_0_n3,
         Red_ToCheckInst_LFInst_1_LFInst_1_n3,
         Red_ToCheckInst_LFInst_1_LFInst_2_n3,
         Red_ToCheckInst_LFInst_2_LFInst_0_n3,
         Red_ToCheckInst_LFInst_2_LFInst_1_n3,
         Red_ToCheckInst_LFInst_2_LFInst_2_n3,
         Red_ToCheckInst_LFInst_3_LFInst_0_n3,
         Red_ToCheckInst_LFInst_3_LFInst_1_n3,
         Red_ToCheckInst_LFInst_3_LFInst_2_n3,
         Red_ToCheckInst_LFInst_4_LFInst_0_n3,
         Red_ToCheckInst_LFInst_4_LFInst_1_n3,
         Red_ToCheckInst_LFInst_4_LFInst_2_n3,
         Red_ToCheckInst_LFInst_5_LFInst_0_n3,
         Red_ToCheckInst_LFInst_5_LFInst_1_n3,
         Red_ToCheckInst_LFInst_5_LFInst_2_n3,
         Red_ToCheckInst_LFInst_6_LFInst_0_n3,
         Red_ToCheckInst_LFInst_6_LFInst_1_n3,
         Red_ToCheckInst_LFInst_6_LFInst_2_n3,
         Red_ToCheckInst_LFInst_7_LFInst_0_n3,
         Red_ToCheckInst_LFInst_7_LFInst_1_n3,
         Red_ToCheckInst_LFInst_7_LFInst_2_n3,
         Red_ToCheckInst_LFInst_8_LFInst_0_n3,
         Red_ToCheckInst_LFInst_8_LFInst_1_n3,
         Red_ToCheckInst_LFInst_8_LFInst_2_n3,
         Red_ToCheckInst_LFInst_9_LFInst_0_n3,
         Red_ToCheckInst_LFInst_9_LFInst_1_n3,
         Red_ToCheckInst_LFInst_9_LFInst_2_n3,
         Red_ToCheckInst_LFInst_10_LFInst_0_n3,
         Red_ToCheckInst_LFInst_10_LFInst_1_n3,
         Red_ToCheckInst_LFInst_10_LFInst_2_n3,
         Red_ToCheckInst_LFInst_11_LFInst_0_n3,
         Red_ToCheckInst_LFInst_11_LFInst_1_n3,
         Red_ToCheckInst_LFInst_11_LFInst_2_n3,
         Red_ToCheckInst_LFInst_12_LFInst_0_n3,
         Red_ToCheckInst_LFInst_12_LFInst_1_n3,
         Red_ToCheckInst_LFInst_12_LFInst_2_n3,
         Red_ToCheckInst_LFInst_13_LFInst_0_n3,
         Red_ToCheckInst_LFInst_13_LFInst_1_n3,
         Red_ToCheckInst_LFInst_13_LFInst_2_n3,
         Red_ToCheckInst_LFInst_14_LFInst_0_n3,
         Red_ToCheckInst_LFInst_14_LFInst_1_n3,
         Red_ToCheckInst_LFInst_14_LFInst_2_n3,
         Red_ToCheckInst_LFInst_15_LFInst_0_n3,
         Red_ToCheckInst_LFInst_15_LFInst_1_n3,
         Red_ToCheckInst_LFInst_15_LFInst_2_n3,
         Red_ToCheckInst_LFInst_16_LFInst_0_n3,
         Red_ToCheckInst_LFInst_16_LFInst_1_n3,
         Red_ToCheckInst_LFInst_16_LFInst_2_n3,
         Red_ToCheckInst_LFInst_17_LFInst_0_n3,
         Red_ToCheckInst_LFInst_17_LFInst_1_n3,
         Red_ToCheckInst_LFInst_17_LFInst_2_n3,
         Red_ToCheckInst_LFInst_18_LFInst_0_n3,
         Red_ToCheckInst_LFInst_18_LFInst_1_n3,
         Red_ToCheckInst_LFInst_18_LFInst_2_n3,
         Red_ToCheckInst_LFInst_19_LFInst_0_n3,
         Red_ToCheckInst_LFInst_19_LFInst_1_n3,
         Red_ToCheckInst_LFInst_19_LFInst_2_n3,
         Red_ToCheckInst_LFInst_20_LFInst_0_n3,
         Red_ToCheckInst_LFInst_20_LFInst_1_n3,
         Red_ToCheckInst_LFInst_20_LFInst_2_n3,
         Red_ToCheckInst_LFInst_21_LFInst_0_n3,
         Red_ToCheckInst_LFInst_21_LFInst_1_n3,
         Red_ToCheckInst_LFInst_21_LFInst_2_n3,
         Red_ToCheckInst_LFInst_22_LFInst_0_n3,
         Red_ToCheckInst_LFInst_22_LFInst_1_n3,
         Red_ToCheckInst_LFInst_22_LFInst_2_n3,
         Red_ToCheckInst_LFInst_23_LFInst_0_n3,
         Red_ToCheckInst_LFInst_23_LFInst_1_n3,
         Red_ToCheckInst_LFInst_23_LFInst_2_n3,
         Red_ToCheckInst_LFInst_24_LFInst_0_n3,
         Red_ToCheckInst_LFInst_24_LFInst_1_n3,
         Red_ToCheckInst_LFInst_24_LFInst_2_n3,
         Red_ToCheckInst_LFInst_25_LFInst_0_n3,
         Red_ToCheckInst_LFInst_25_LFInst_1_n3,
         Red_ToCheckInst_LFInst_25_LFInst_2_n3,
         Red_ToCheckInst_LFInst_26_LFInst_0_n3,
         Red_ToCheckInst_LFInst_26_LFInst_1_n3,
         Red_ToCheckInst_LFInst_26_LFInst_2_n3,
         Red_ToCheckInst_LFInst_27_LFInst_0_n3,
         Red_ToCheckInst_LFInst_27_LFInst_1_n3,
         Red_ToCheckInst_LFInst_27_LFInst_2_n3,
         Red_ToCheckInst_LFInst_28_LFInst_0_n3,
         Red_ToCheckInst_LFInst_28_LFInst_1_n3,
         Red_ToCheckInst_LFInst_28_LFInst_2_n3,
         Red_ToCheckInst_LFInst_29_LFInst_0_n3,
         Red_ToCheckInst_LFInst_29_LFInst_1_n3,
         Red_ToCheckInst_LFInst_29_LFInst_2_n3,
         Red_ToCheckInst_LFInst_30_LFInst_0_n3,
         Red_ToCheckInst_LFInst_30_LFInst_1_n3,
         Red_ToCheckInst_LFInst_30_LFInst_2_n3,
         Red_ToCheckInst_LFInst_31_LFInst_0_n3,
         Red_ToCheckInst_LFInst_31_LFInst_1_n3,
         Red_ToCheckInst_LFInst_31_LFInst_2_n3,
         Red_ToCheckInst_LFInst_32_LFInst_0_n3,
         Red_ToCheckInst_LFInst_32_LFInst_1_n3,
         Red_ToCheckInst_LFInst_32_LFInst_2_n3,
         Red_ToCheckInst_LFInst_33_LFInst_0_n3,
         Red_ToCheckInst_LFInst_33_LFInst_1_n3,
         Red_ToCheckInst_LFInst_33_LFInst_2_n3,
         Red_ToCheckInst_LFInst_34_LFInst_0_n3,
         Red_ToCheckInst_LFInst_34_LFInst_1_n3,
         Red_ToCheckInst_LFInst_34_LFInst_2_n3,
         Red_ToCheckInst_LFInst_35_LFInst_0_n3,
         Red_ToCheckInst_LFInst_35_LFInst_1_n3,
         Red_ToCheckInst_LFInst_35_LFInst_2_n3,
         Red_ToCheckInst_LFInst_36_LFInst_0_n3,
         Red_ToCheckInst_LFInst_36_LFInst_1_n3,
         Red_ToCheckInst_LFInst_36_LFInst_2_n3,
         Red_ToCheckInst_LFInst_37_LFInst_0_n3,
         Red_ToCheckInst_LFInst_37_LFInst_1_n3,
         Red_ToCheckInst_LFInst_37_LFInst_2_n3,
         Red_ToCheckInst_LFInst_38_LFInst_0_n3,
         Red_ToCheckInst_LFInst_38_LFInst_1_n3,
         Red_ToCheckInst_LFInst_38_LFInst_2_n3,
         Red_ToCheckInst_LFInst_39_LFInst_0_n3,
         Red_ToCheckInst_LFInst_39_LFInst_1_n3,
         Red_ToCheckInst_LFInst_39_LFInst_2_n3,
         Red_ToCheckInst_LFInst_40_LFInst_0_n3,
         Red_ToCheckInst_LFInst_40_LFInst_1_n3,
         Red_ToCheckInst_LFInst_40_LFInst_2_n3,
         Red_ToCheckInst_LFInst_41_LFInst_0_n3,
         Red_ToCheckInst_LFInst_41_LFInst_1_n3,
         Red_ToCheckInst_LFInst_41_LFInst_2_n3,
         Red_ToCheckInst_LFInst_42_LFInst_0_n3,
         Red_ToCheckInst_LFInst_42_LFInst_1_n3,
         Red_ToCheckInst_LFInst_42_LFInst_2_n3,
         Red_ToCheckInst_LFInst_43_LFInst_0_n3,
         Red_ToCheckInst_LFInst_43_LFInst_1_n3,
         Red_ToCheckInst_LFInst_43_LFInst_2_n3,
         Red_ToCheckInst_LFInst_44_LFInst_0_n3,
         Red_ToCheckInst_LFInst_44_LFInst_1_n3,
         Red_ToCheckInst_LFInst_44_LFInst_2_n3,
         Red_ToCheckInst_LFInst_45_LFInst_0_n3,
         Red_ToCheckInst_LFInst_45_LFInst_1_n3,
         Red_ToCheckInst_LFInst_45_LFInst_2_n3,
         Red_ToCheckInst_LFInst_46_LFInst_0_n3,
         Red_ToCheckInst_LFInst_46_LFInst_1_n3,
         Red_ToCheckInst_LFInst_46_LFInst_2_n3,
         Red_ToCheckInst_LFInst_47_LFInst_0_n3,
         Red_ToCheckInst_LFInst_47_LFInst_1_n3,
         Red_ToCheckInst_LFInst_47_LFInst_2_n3,
         Red_ToCheckInst_LFInst_48_LFInst_0_n3,
         Red_ToCheckInst_LFInst_48_LFInst_1_n3,
         Red_ToCheckInst_LFInst_48_LFInst_2_n3,
         Red_ToCheckInst_LFInst_49_LFInst_0_n3,
         Red_ToCheckInst_LFInst_49_LFInst_1_n3,
         Red_ToCheckInst_LFInst_49_LFInst_2_n3,
         Red_ToCheckInst_LFInst_50_LFInst_0_n3,
         Red_ToCheckInst_LFInst_50_LFInst_1_n3,
         Red_ToCheckInst_LFInst_50_LFInst_2_n3,
         Red_ToCheckInst_LFInst_51_LFInst_0_n3,
         Red_ToCheckInst_LFInst_51_LFInst_1_n3,
         Red_ToCheckInst_LFInst_51_LFInst_2_n3,
         Red_ToCheckInst_LFInst_52_LFInst_0_n3,
         Red_ToCheckInst_LFInst_52_LFInst_1_n3,
         Red_ToCheckInst_LFInst_52_LFInst_2_n3,
         Red_ToCheckInst_LFInst_53_LFInst_0_n3,
         Red_ToCheckInst_LFInst_53_LFInst_1_n3,
         Red_ToCheckInst_LFInst_53_LFInst_2_n3,
         Red_ToCheckInst_LFInst_54_LFInst_0_n3,
         Red_ToCheckInst_LFInst_54_LFInst_1_n3,
         Red_ToCheckInst_LFInst_54_LFInst_2_n3,
         Red_ToCheckInst_LFInst_55_LFInst_0_n3,
         Red_ToCheckInst_LFInst_55_LFInst_1_n3,
         Red_ToCheckInst_LFInst_55_LFInst_2_n3,
         Red_ToCheckInst_LFInst_56_LFInst_0_n3,
         Red_ToCheckInst_LFInst_56_LFInst_1_n3,
         Red_ToCheckInst_LFInst_56_LFInst_2_n3,
         Red_ToCheckInst_LFInst_57_LFInst_0_n3,
         Red_ToCheckInst_LFInst_57_LFInst_1_n3,
         Red_ToCheckInst_LFInst_57_LFInst_2_n3,
         Red_ToCheckInst_LFInst_58_LFInst_0_n3,
         Red_ToCheckInst_LFInst_58_LFInst_1_n3,
         Red_ToCheckInst_LFInst_58_LFInst_2_n3,
         Red_ToCheckInst_LFInst_59_LFInst_0_n3,
         Red_ToCheckInst_LFInst_59_LFInst_1_n3,
         Red_ToCheckInst_LFInst_59_LFInst_2_n3,
         Red_ToCheckInst_LFInst_60_LFInst_0_n3,
         Red_ToCheckInst_LFInst_60_LFInst_1_n3,
         Red_ToCheckInst_LFInst_60_LFInst_2_n3,
         Red_ToCheckInst_LFInst_61_LFInst_0_n3,
         Red_ToCheckInst_LFInst_61_LFInst_1_n3,
         Red_ToCheckInst_LFInst_61_LFInst_2_n3,
         Red_ToCheckInst_LFInst_62_LFInst_0_n3,
         Red_ToCheckInst_LFInst_62_LFInst_1_n3,
         Red_ToCheckInst_LFInst_62_LFInst_2_n3,
         Red_ToCheckInst_LFInst_63_LFInst_0_n3,
         Red_ToCheckInst_LFInst_63_LFInst_1_n3,
         Red_ToCheckInst_LFInst_63_LFInst_2_n3,
         Red_ToCheckInst_LFInst_64_LFInst_0_n3,
         Red_ToCheckInst_LFInst_64_LFInst_1_n3,
         Red_ToCheckInst_LFInst_64_LFInst_2_n3,
         Red_ToCheckInst_LFInst_65_LFInst_0_n3,
         Red_ToCheckInst_LFInst_65_LFInst_1_n3,
         Red_ToCheckInst_LFInst_65_LFInst_2_n3,
         Red_ToCheckInst_LFInst_66_LFInst_0_n3,
         Red_ToCheckInst_LFInst_66_LFInst_1_n3,
         Red_ToCheckInst_LFInst_66_LFInst_2_n3,
         Red_ToCheckInst_LFInst_67_LFInst_0_n3,
         Red_ToCheckInst_LFInst_67_LFInst_1_n3,
         Red_ToCheckInst_LFInst_67_LFInst_2_n3,
         Red_ToCheckInst_LFInst_68_LFInst_0_n3,
         Red_ToCheckInst_LFInst_68_LFInst_1_n3,
         Red_ToCheckInst_LFInst_68_LFInst_2_n3,
         Red_ToCheckInst_LFInst_69_LFInst_0_n3,
         Red_ToCheckInst_LFInst_69_LFInst_1_n3,
         Red_ToCheckInst_LFInst_69_LFInst_2_n3,
         Red_ToCheckInst_LFInst_70_LFInst_0_n3,
         Red_ToCheckInst_LFInst_70_LFInst_1_n3,
         Red_ToCheckInst_LFInst_70_LFInst_2_n3,
         Red_ToCheckInst_LFInst_71_LFInst_0_n3,
         Red_ToCheckInst_LFInst_71_LFInst_1_n3,
         Red_ToCheckInst_LFInst_71_LFInst_2_n3,
         Red_ToCheckInst_LFInst_72_LFInst_0_n3,
         Red_ToCheckInst_LFInst_72_LFInst_1_n3,
         Red_ToCheckInst_LFInst_72_LFInst_2_n3,
         Red_ToCheckInst_LFInst_73_LFInst_0_n3,
         Red_ToCheckInst_LFInst_73_LFInst_1_n3,
         Red_ToCheckInst_LFInst_73_LFInst_2_n3,
         Red_ToCheckInst_LFInst_74_LFInst_0_n3,
         Red_ToCheckInst_LFInst_74_LFInst_1_n3,
         Red_ToCheckInst_LFInst_74_LFInst_2_n3,
         Red_ToCheckInst_LFInst_75_LFInst_0_n3,
         Red_ToCheckInst_LFInst_75_LFInst_1_n3,
         Red_ToCheckInst_LFInst_75_LFInst_2_n3,
         Red_ToCheckInst_LFInst_76_LFInst_0_n3,
         Red_ToCheckInst_LFInst_76_LFInst_1_n3,
         Red_ToCheckInst_LFInst_76_LFInst_2_n3,
         Red_ToCheckInst_LFInst_77_LFInst_0_n3,
         Red_ToCheckInst_LFInst_77_LFInst_1_n3,
         Red_ToCheckInst_LFInst_77_LFInst_2_n3,
         Red_ToCheckInst_LFInst_78_LFInst_0_n3,
         Red_ToCheckInst_LFInst_78_LFInst_1_n3,
         Red_ToCheckInst_LFInst_78_LFInst_2_n3,
         Red_ToCheckInst_LFInst_79_LFInst_0_n3,
         Red_ToCheckInst_LFInst_79_LFInst_1_n3,
         Red_ToCheckInst_LFInst_79_LFInst_2_n3,
         Red_ToCheckInst_LFInst_80_LFInst_0_n3,
         Red_ToCheckInst_LFInst_80_LFInst_1_n3,
         Red_ToCheckInst_LFInst_80_LFInst_2_n3,
         Red_ToCheckInst_LFInst_81_LFInst_0_n3,
         Red_ToCheckInst_LFInst_81_LFInst_1_n3,
         Red_ToCheckInst_LFInst_81_LFInst_2_n3,
         Red_ToCheckInst_LFInst_82_LFInst_0_n3,
         Red_ToCheckInst_LFInst_82_LFInst_1_n3,
         Red_ToCheckInst_LFInst_82_LFInst_2_n3,
         Red_ToCheckInst_LFInst_83_LFInst_0_n3,
         Red_ToCheckInst_LFInst_83_LFInst_1_n3,
         Red_ToCheckInst_LFInst_83_LFInst_2_n3,
         Red_ToCheckInst_LFInst_84_LFInst_0_n3,
         Red_ToCheckInst_LFInst_84_LFInst_1_n3,
         Red_ToCheckInst_LFInst_84_LFInst_2_n3,
         Red_ToCheckInst_LFInst_85_LFInst_0_n3,
         Red_ToCheckInst_LFInst_85_LFInst_1_n3,
         Red_ToCheckInst_LFInst_85_LFInst_2_n3,
         Red_ToCheckInst_LFInst_86_LFInst_0_n3,
         Red_ToCheckInst_LFInst_86_LFInst_1_n3,
         Red_ToCheckInst_LFInst_86_LFInst_2_n3,
         Red_ToCheckInst_LFInst_87_LFInst_0_n3,
         Red_ToCheckInst_LFInst_87_LFInst_1_n3,
         Red_ToCheckInst_LFInst_87_LFInst_2_n3,
         Red_ToCheckInst_LFInst_88_LFInst_0_n3,
         Red_ToCheckInst_LFInst_88_LFInst_1_n3,
         Red_ToCheckInst_LFInst_88_LFInst_2_n3,
         Red_ToCheckInst_LFInst_89_LFInst_0_n3,
         Red_ToCheckInst_LFInst_89_LFInst_1_n3,
         Red_ToCheckInst_LFInst_89_LFInst_2_n3,
         Red_ToCheckInst_LFInst_90_LFInst_0_n3,
         Red_ToCheckInst_LFInst_90_LFInst_1_n3,
         Red_ToCheckInst_LFInst_90_LFInst_2_n3,
         Red_ToCheckInst_LFInst_91_LFInst_0_n3,
         Red_ToCheckInst_LFInst_91_LFInst_1_n3,
         Red_ToCheckInst_LFInst_91_LFInst_2_n3,
         Red_ToCheckInst_LFInst_92_LFInst_0_n3,
         Red_ToCheckInst_LFInst_92_LFInst_1_n3,
         Red_ToCheckInst_LFInst_92_LFInst_2_n3,
         Red_ToCheckInst_LFInst_93_LFInst_0_n3,
         Red_ToCheckInst_LFInst_93_LFInst_1_n3,
         Red_ToCheckInst_LFInst_93_LFInst_2_n3,
         Red_ToCheckInst_LFInst_94_LFInst_0_n3,
         Red_ToCheckInst_LFInst_94_LFInst_1_n3,
         Red_ToCheckInst_LFInst_94_LFInst_2_n3,
         Red_ToCheckInst_LFInst_95_LFInst_0_n3,
         Red_ToCheckInst_LFInst_95_LFInst_1_n3,
         Red_ToCheckInst_LFInst_95_LFInst_2_n3, Check1_CheckInst_0_n190,
         Check1_CheckInst_0_n189, Check1_CheckInst_0_n188,
         Check1_CheckInst_0_n187, Check1_CheckInst_0_n186,
         Check1_CheckInst_0_n185, Check1_CheckInst_0_n184,
         Check1_CheckInst_0_n183, Check1_CheckInst_0_n182,
         Check1_CheckInst_0_n181, Check1_CheckInst_0_n180,
         Check1_CheckInst_0_n179, Check1_CheckInst_0_n178,
         Check1_CheckInst_0_n177, Check1_CheckInst_0_n176,
         Check1_CheckInst_0_n175, Check1_CheckInst_0_n174,
         Check1_CheckInst_0_n173, Check1_CheckInst_0_n172,
         Check1_CheckInst_0_n171, Check1_CheckInst_0_n170,
         Check1_CheckInst_0_n169, Check1_CheckInst_0_n168,
         Check1_CheckInst_0_n167, Check1_CheckInst_0_n166,
         Check1_CheckInst_0_n165, Check1_CheckInst_0_n164,
         Check1_CheckInst_0_n163, Check1_CheckInst_0_n162,
         Check1_CheckInst_0_n161, Check1_CheckInst_0_n160,
         Check1_CheckInst_0_n159, Check1_CheckInst_0_n158,
         Check1_CheckInst_0_n157, Check1_CheckInst_0_n156,
         Check1_CheckInst_0_n155, Check1_CheckInst_0_n154,
         Check1_CheckInst_0_n153, Check1_CheckInst_0_n152,
         Check1_CheckInst_0_n151, Check1_CheckInst_0_n150,
         Check1_CheckInst_0_n149, Check1_CheckInst_0_n148,
         Check1_CheckInst_0_n147, Check1_CheckInst_0_n146,
         Check1_CheckInst_0_n145, Check1_CheckInst_0_n144,
         Check1_CheckInst_0_n143, Check1_CheckInst_0_n142,
         Check1_CheckInst_0_n141, Check1_CheckInst_0_n140,
         Check1_CheckInst_0_n139, Check1_CheckInst_0_n138,
         Check1_CheckInst_0_n137, Check1_CheckInst_0_n136,
         Check1_CheckInst_0_n135, Check1_CheckInst_0_n134,
         Check1_CheckInst_0_n133, Check1_CheckInst_0_n132,
         Check1_CheckInst_0_n131, Check1_CheckInst_0_n130,
         Check1_CheckInst_0_n129, Check1_CheckInst_0_n128,
         Check1_CheckInst_0_n127, Check1_CheckInst_0_n126,
         Check1_CheckInst_0_n125, Check1_CheckInst_0_n124,
         Check1_CheckInst_0_n123, Check1_CheckInst_0_n122,
         Check1_CheckInst_0_n121, Check1_CheckInst_0_n120,
         Check1_CheckInst_0_n119, Check1_CheckInst_0_n118,
         Check1_CheckInst_0_n117, Check1_CheckInst_0_n116,
         Check1_CheckInst_0_n115, Check1_CheckInst_0_n114,
         Check1_CheckInst_0_n113, Check1_CheckInst_0_n112,
         Check1_CheckInst_0_n111, Check1_CheckInst_0_n110,
         Check1_CheckInst_0_n109, Check1_CheckInst_0_n108,
         Check1_CheckInst_0_n107, Check1_CheckInst_0_n106,
         Check1_CheckInst_0_n105, Check1_CheckInst_0_n104,
         Check1_CheckInst_0_n103, Check1_CheckInst_0_n102,
         Check1_CheckInst_0_n101, Check1_CheckInst_0_n100,
         Check1_CheckInst_0_n99, Check1_CheckInst_0_n98,
         Check1_CheckInst_0_n97, Check1_CheckInst_0_n96,
         Check1_CheckInst_0_n95, Check1_CheckInst_0_n94,
         Check1_CheckInst_0_n93, Check1_CheckInst_0_n92,
         Check1_CheckInst_0_n91, Check1_CheckInst_0_n90,
         Check1_CheckInst_0_n89, Check1_CheckInst_0_n88,
         Check1_CheckInst_0_n87, Check1_CheckInst_0_n86,
         Check1_CheckInst_0_n85, Check1_CheckInst_0_n84,
         Check1_CheckInst_0_n83, Check1_CheckInst_0_n82,
         Check1_CheckInst_0_n81, Check1_CheckInst_0_n80,
         Check1_CheckInst_0_n79, Check1_CheckInst_0_n78,
         Check1_CheckInst_0_n77, Check1_CheckInst_0_n76,
         Check1_CheckInst_0_n75, Check1_CheckInst_0_n74,
         Check1_CheckInst_0_n73, Check1_CheckInst_0_n72,
         Check1_CheckInst_0_n71, Check1_CheckInst_0_n70,
         Check1_CheckInst_0_n69, Check1_CheckInst_0_n68,
         Check1_CheckInst_0_n67, Check1_CheckInst_0_n66,
         Check1_CheckInst_0_n65, Check1_CheckInst_0_n64,
         Check1_CheckInst_0_n63, Check1_CheckInst_0_n62,
         Check1_CheckInst_0_n61, Check1_CheckInst_0_n60,
         Check1_CheckInst_0_n59, Check1_CheckInst_0_n58,
         Check1_CheckInst_0_n57, Check1_CheckInst_0_n56,
         Check1_CheckInst_0_n55, Check1_CheckInst_0_n54,
         Check1_CheckInst_0_n53, Check1_CheckInst_0_n52,
         Check1_CheckInst_0_n51, Check1_CheckInst_0_n50,
         Check1_CheckInst_0_n49, Check1_CheckInst_0_n48,
         Check1_CheckInst_0_n47, Check1_CheckInst_0_n46,
         Check1_CheckInst_0_n45, Check1_CheckInst_0_n44,
         Check1_CheckInst_0_n43, Check1_CheckInst_0_n42,
         Check1_CheckInst_0_n41, Check1_CheckInst_0_n40,
         Check1_CheckInst_0_n39, Check1_CheckInst_0_n38,
         Check1_CheckInst_0_n37, Check1_CheckInst_0_n36,
         Check1_CheckInst_0_n35, Check1_CheckInst_0_n34,
         Check1_CheckInst_0_n33, Check1_CheckInst_0_n32,
         Check1_CheckInst_0_n31, Check1_CheckInst_0_n30,
         Check1_CheckInst_0_n29, Check1_CheckInst_0_n28,
         Check1_CheckInst_0_n27, Check1_CheckInst_0_n26,
         Check1_CheckInst_0_n25, Check1_CheckInst_0_n24,
         Check1_CheckInst_0_n23, Check1_CheckInst_0_n22,
         Check1_CheckInst_0_n21, Check1_CheckInst_0_n20,
         Check1_CheckInst_0_n19, Check1_CheckInst_0_n18,
         Check1_CheckInst_0_n17, Check1_CheckInst_0_n16,
         Check1_CheckInst_0_n15, Check1_CheckInst_0_n14,
         Check1_CheckInst_0_n13, Check1_CheckInst_0_n12,
         Check1_CheckInst_0_n11, Check1_CheckInst_0_n10, Check1_CheckInst_0_n9,
         Check1_CheckInst_0_n8, Check1_CheckInst_0_n7, Check1_CheckInst_0_n6,
         Check1_CheckInst_0_n5, Check1_CheckInst_0_n4, Check1_CheckInst_0_n3,
         Check1_CheckInst_0_n2, Check1_CheckInst_0_n1, Check1_CheckInst_1_n192,
         Check1_CheckInst_1_n191, Check1_CheckInst_1_n190,
         Check1_CheckInst_1_n189, Check1_CheckInst_1_n188,
         Check1_CheckInst_1_n187, Check1_CheckInst_1_n186,
         Check1_CheckInst_1_n185, Check1_CheckInst_1_n184,
         Check1_CheckInst_1_n183, Check1_CheckInst_1_n182,
         Check1_CheckInst_1_n181, Check1_CheckInst_1_n180,
         Check1_CheckInst_1_n179, Check1_CheckInst_1_n178,
         Check1_CheckInst_1_n177, Check1_CheckInst_1_n176,
         Check1_CheckInst_1_n175, Check1_CheckInst_1_n174,
         Check1_CheckInst_1_n173, Check1_CheckInst_1_n172,
         Check1_CheckInst_1_n171, Check1_CheckInst_1_n170,
         Check1_CheckInst_1_n169, Check1_CheckInst_1_n168,
         Check1_CheckInst_1_n167, Check1_CheckInst_1_n166,
         Check1_CheckInst_1_n165, Check1_CheckInst_1_n164,
         Check1_CheckInst_1_n163, Check1_CheckInst_1_n162,
         Check1_CheckInst_1_n161, Check1_CheckInst_1_n160,
         Check1_CheckInst_1_n159, Check1_CheckInst_1_n158,
         Check1_CheckInst_1_n157, Check1_CheckInst_1_n156,
         Check1_CheckInst_1_n155, Check1_CheckInst_1_n154,
         Check1_CheckInst_1_n153, Check1_CheckInst_1_n152,
         Check1_CheckInst_1_n151, Check1_CheckInst_1_n150,
         Check1_CheckInst_1_n149, Check1_CheckInst_1_n148,
         Check1_CheckInst_1_n147, Check1_CheckInst_1_n146,
         Check1_CheckInst_1_n145, Check1_CheckInst_1_n144,
         Check1_CheckInst_1_n143, Check1_CheckInst_1_n142,
         Check1_CheckInst_1_n141, Check1_CheckInst_1_n140,
         Check1_CheckInst_1_n139, Check1_CheckInst_1_n138,
         Check1_CheckInst_1_n137, Check1_CheckInst_1_n136,
         Check1_CheckInst_1_n135, Check1_CheckInst_1_n134,
         Check1_CheckInst_1_n133, Check1_CheckInst_1_n132,
         Check1_CheckInst_1_n131, Check1_CheckInst_1_n130,
         Check1_CheckInst_1_n129, Check1_CheckInst_1_n128,
         Check1_CheckInst_1_n127, Check1_CheckInst_1_n126,
         Check1_CheckInst_1_n125, Check1_CheckInst_1_n124,
         Check1_CheckInst_1_n123, Check1_CheckInst_1_n122,
         Check1_CheckInst_1_n121, Check1_CheckInst_1_n120,
         Check1_CheckInst_1_n119, Check1_CheckInst_1_n118,
         Check1_CheckInst_1_n117, Check1_CheckInst_1_n116,
         Check1_CheckInst_1_n115, Check1_CheckInst_1_n114,
         Check1_CheckInst_1_n113, Check1_CheckInst_1_n112,
         Check1_CheckInst_1_n111, Check1_CheckInst_1_n110,
         Check1_CheckInst_1_n109, Check1_CheckInst_1_n108,
         Check1_CheckInst_1_n107, Check1_CheckInst_1_n106,
         Check1_CheckInst_1_n105, Check1_CheckInst_1_n104,
         Check1_CheckInst_1_n103, Check1_CheckInst_1_n102,
         Check1_CheckInst_1_n101, Check1_CheckInst_1_n100,
         Check1_CheckInst_1_n99, Check1_CheckInst_1_n98,
         Check1_CheckInst_1_n97, Check1_CheckInst_1_n96,
         Check1_CheckInst_1_n95, Check1_CheckInst_1_n94,
         Check1_CheckInst_1_n93, Check1_CheckInst_1_n92,
         Check1_CheckInst_1_n91, Check1_CheckInst_1_n90,
         Check1_CheckInst_1_n89, Check1_CheckInst_1_n88,
         Check1_CheckInst_1_n87, Check1_CheckInst_1_n86,
         Check1_CheckInst_1_n85, Check1_CheckInst_1_n84,
         Check1_CheckInst_1_n83, Check1_CheckInst_1_n82,
         Check1_CheckInst_1_n81, Check1_CheckInst_1_n80,
         Check1_CheckInst_1_n79, Check1_CheckInst_1_n78,
         Check1_CheckInst_1_n77, Check1_CheckInst_1_n76,
         Check1_CheckInst_1_n75, Check1_CheckInst_1_n74,
         Check1_CheckInst_1_n73, Check1_CheckInst_1_n72,
         Check1_CheckInst_1_n71, Check1_CheckInst_1_n70,
         Check1_CheckInst_1_n69, Check1_CheckInst_1_n68,
         Check1_CheckInst_1_n67, Check1_CheckInst_1_n66,
         Check1_CheckInst_1_n65, Check1_CheckInst_1_n64,
         Check1_CheckInst_1_n63, Check1_CheckInst_1_n62,
         Check1_CheckInst_1_n61, Check1_CheckInst_1_n60,
         Check1_CheckInst_1_n59, Check1_CheckInst_1_n58,
         Check1_CheckInst_1_n57, Check1_CheckInst_1_n56,
         Check1_CheckInst_1_n55, Check1_CheckInst_1_n54,
         Check1_CheckInst_1_n53, Check1_CheckInst_1_n52,
         Check1_CheckInst_1_n51, Check1_CheckInst_1_n50,
         Check1_CheckInst_1_n49, Check1_CheckInst_1_n48,
         Check1_CheckInst_1_n47, Check1_CheckInst_1_n46,
         Check1_CheckInst_1_n45, Check1_CheckInst_1_n44,
         Check1_CheckInst_1_n43, Check1_CheckInst_1_n42,
         Check1_CheckInst_1_n41, Check1_CheckInst_1_n40,
         Check1_CheckInst_1_n39, Check1_CheckInst_1_n38,
         Check1_CheckInst_1_n37, Check1_CheckInst_1_n36,
         Check1_CheckInst_1_n35, Check1_CheckInst_1_n34,
         Check1_CheckInst_1_n33, Check1_CheckInst_1_n32,
         Check1_CheckInst_1_n31, Check1_CheckInst_1_n30,
         Check1_CheckInst_1_n29, Check1_CheckInst_1_n28,
         Check1_CheckInst_1_n27, Check1_CheckInst_1_n26,
         Check1_CheckInst_1_n25, Check1_CheckInst_1_n24,
         Check1_CheckInst_1_n23, Check1_CheckInst_1_n22,
         Check1_CheckInst_1_n21, Check1_CheckInst_1_n20,
         Check1_CheckInst_1_n19, Check1_CheckInst_1_n18,
         Check1_CheckInst_1_n17, Check1_CheckInst_1_n16,
         Check1_CheckInst_1_n15, Check1_CheckInst_1_n14,
         Check1_CheckInst_1_n13, Check1_CheckInst_1_n12,
         Check1_CheckInst_1_n11, Check1_CheckInst_1_n10, Check1_CheckInst_1_n9,
         Check1_CheckInst_1_n8, Check1_CheckInst_1_n7, Check1_CheckInst_1_n6,
         Check1_CheckInst_1_n5, Check1_CheckInst_1_n4, Check1_CheckInst_1_n3,
         Check1_CheckInst_2_n192, Check1_CheckInst_2_n191,
         Check1_CheckInst_2_n190, Check1_CheckInst_2_n189,
         Check1_CheckInst_2_n188, Check1_CheckInst_2_n187,
         Check1_CheckInst_2_n186, Check1_CheckInst_2_n185,
         Check1_CheckInst_2_n184, Check1_CheckInst_2_n183,
         Check1_CheckInst_2_n182, Check1_CheckInst_2_n181,
         Check1_CheckInst_2_n180, Check1_CheckInst_2_n179,
         Check1_CheckInst_2_n178, Check1_CheckInst_2_n177,
         Check1_CheckInst_2_n176, Check1_CheckInst_2_n175,
         Check1_CheckInst_2_n174, Check1_CheckInst_2_n173,
         Check1_CheckInst_2_n172, Check1_CheckInst_2_n171,
         Check1_CheckInst_2_n170, Check1_CheckInst_2_n169,
         Check1_CheckInst_2_n168, Check1_CheckInst_2_n167,
         Check1_CheckInst_2_n166, Check1_CheckInst_2_n165,
         Check1_CheckInst_2_n164, Check1_CheckInst_2_n163,
         Check1_CheckInst_2_n162, Check1_CheckInst_2_n161,
         Check1_CheckInst_2_n160, Check1_CheckInst_2_n159,
         Check1_CheckInst_2_n158, Check1_CheckInst_2_n157,
         Check1_CheckInst_2_n156, Check1_CheckInst_2_n155,
         Check1_CheckInst_2_n154, Check1_CheckInst_2_n153,
         Check1_CheckInst_2_n152, Check1_CheckInst_2_n151,
         Check1_CheckInst_2_n150, Check1_CheckInst_2_n149,
         Check1_CheckInst_2_n148, Check1_CheckInst_2_n147,
         Check1_CheckInst_2_n146, Check1_CheckInst_2_n145,
         Check1_CheckInst_2_n144, Check1_CheckInst_2_n143,
         Check1_CheckInst_2_n142, Check1_CheckInst_2_n141,
         Check1_CheckInst_2_n140, Check1_CheckInst_2_n139,
         Check1_CheckInst_2_n138, Check1_CheckInst_2_n137,
         Check1_CheckInst_2_n136, Check1_CheckInst_2_n135,
         Check1_CheckInst_2_n134, Check1_CheckInst_2_n133,
         Check1_CheckInst_2_n132, Check1_CheckInst_2_n131,
         Check1_CheckInst_2_n130, Check1_CheckInst_2_n129,
         Check1_CheckInst_2_n128, Check1_CheckInst_2_n127,
         Check1_CheckInst_2_n126, Check1_CheckInst_2_n125,
         Check1_CheckInst_2_n124, Check1_CheckInst_2_n123,
         Check1_CheckInst_2_n122, Check1_CheckInst_2_n121,
         Check1_CheckInst_2_n120, Check1_CheckInst_2_n119,
         Check1_CheckInst_2_n118, Check1_CheckInst_2_n117,
         Check1_CheckInst_2_n116, Check1_CheckInst_2_n115,
         Check1_CheckInst_2_n114, Check1_CheckInst_2_n113,
         Check1_CheckInst_2_n112, Check1_CheckInst_2_n111,
         Check1_CheckInst_2_n110, Check1_CheckInst_2_n109,
         Check1_CheckInst_2_n108, Check1_CheckInst_2_n107,
         Check1_CheckInst_2_n106, Check1_CheckInst_2_n105,
         Check1_CheckInst_2_n104, Check1_CheckInst_2_n103,
         Check1_CheckInst_2_n102, Check1_CheckInst_2_n101,
         Check1_CheckInst_2_n100, Check1_CheckInst_2_n99,
         Check1_CheckInst_2_n98, Check1_CheckInst_2_n97,
         Check1_CheckInst_2_n96, Check1_CheckInst_2_n95,
         Check1_CheckInst_2_n94, Check1_CheckInst_2_n93,
         Check1_CheckInst_2_n92, Check1_CheckInst_2_n91,
         Check1_CheckInst_2_n90, Check1_CheckInst_2_n89,
         Check1_CheckInst_2_n88, Check1_CheckInst_2_n87,
         Check1_CheckInst_2_n86, Check1_CheckInst_2_n85,
         Check1_CheckInst_2_n84, Check1_CheckInst_2_n83,
         Check1_CheckInst_2_n82, Check1_CheckInst_2_n81,
         Check1_CheckInst_2_n80, Check1_CheckInst_2_n79,
         Check1_CheckInst_2_n78, Check1_CheckInst_2_n77,
         Check1_CheckInst_2_n76, Check1_CheckInst_2_n75,
         Check1_CheckInst_2_n74, Check1_CheckInst_2_n73,
         Check1_CheckInst_2_n72, Check1_CheckInst_2_n71,
         Check1_CheckInst_2_n70, Check1_CheckInst_2_n69,
         Check1_CheckInst_2_n68, Check1_CheckInst_2_n67,
         Check1_CheckInst_2_n66, Check1_CheckInst_2_n65,
         Check1_CheckInst_2_n64, Check1_CheckInst_2_n63,
         Check1_CheckInst_2_n62, Check1_CheckInst_2_n61,
         Check1_CheckInst_2_n60, Check1_CheckInst_2_n59,
         Check1_CheckInst_2_n58, Check1_CheckInst_2_n57,
         Check1_CheckInst_2_n56, Check1_CheckInst_2_n55,
         Check1_CheckInst_2_n54, Check1_CheckInst_2_n53,
         Check1_CheckInst_2_n52, Check1_CheckInst_2_n51,
         Check1_CheckInst_2_n50, Check1_CheckInst_2_n49,
         Check1_CheckInst_2_n48, Check1_CheckInst_2_n47,
         Check1_CheckInst_2_n46, Check1_CheckInst_2_n45,
         Check1_CheckInst_2_n44, Check1_CheckInst_2_n43,
         Check1_CheckInst_2_n42, Check1_CheckInst_2_n41,
         Check1_CheckInst_2_n40, Check1_CheckInst_2_n39,
         Check1_CheckInst_2_n38, Check1_CheckInst_2_n37,
         Check1_CheckInst_2_n36, Check1_CheckInst_2_n35,
         Check1_CheckInst_2_n34, Check1_CheckInst_2_n33,
         Check1_CheckInst_2_n32, Check1_CheckInst_2_n31,
         Check1_CheckInst_2_n30, Check1_CheckInst_2_n29,
         Check1_CheckInst_2_n28, Check1_CheckInst_2_n27,
         Check1_CheckInst_2_n26, Check1_CheckInst_2_n25,
         Check1_CheckInst_2_n24, Check1_CheckInst_2_n23,
         Check1_CheckInst_2_n22, Check1_CheckInst_2_n21,
         Check1_CheckInst_2_n20, Check1_CheckInst_2_n19,
         Check1_CheckInst_2_n18, Check1_CheckInst_2_n17,
         Check1_CheckInst_2_n16, Check1_CheckInst_2_n15,
         Check1_CheckInst_2_n14, Check1_CheckInst_2_n13,
         Check1_CheckInst_2_n12, Check1_CheckInst_2_n11,
         Check1_CheckInst_2_n10, Check1_CheckInst_2_n9, Check1_CheckInst_2_n8,
         Check1_CheckInst_2_n7, Check1_CheckInst_2_n6, Check1_CheckInst_2_n5,
         Check1_CheckInst_2_n4, Check1_CheckInst_2_n3;
  wire   [63:0] AddRoundKeyOutput;
  wire   [28:16] ShiftRowsOutput;
  wire   [63:0] MC_output;
  wire   [63:0] SubCellInput2;
  wire   [28:16] ShiftRowsOutput2;
  wire   [47:0] Red_Plaintext;
  wire   [47:0] Red_RoundKey;
  wire   [47:0] Red_AddRoundKeyOutput;
  wire   [47:0] Red_ShiftRowsOutput;
  wire   [47:0] Red_MC_output;
  wire   [47:0] Red_SubCellInput2;
  wire   [47:0] Red_ShiftRowsOutput2;
  wire   [47:0] Red_MC_output2;
  wire   [287:0] Red_SignaltoCheck;
  wire   [2:0] Error;
  wire   [3:0] MCInst_MC0_v3_3;
  wire   [3:0] MCInst_MC0_v3_2;
  wire   [3:0] MCInst_MC0_v3_1;
  wire   [3:1] MCInst_MC0_v3_0;
  wire   [3:0] MCInst_MC0_v2_3;
  wire   [3:0] MCInst_MC0_v2_2;
  wire   [3:0] MCInst_MC0_v2_1;
  wire   [3:1] MCInst_MC0_v2_0;
  wire   [3:1] MCInst_MC0_v1_3;
  wire   [3:0] MCInst_MC0_v1_2;
  wire   [3:0] MCInst_MC0_v1_1;
  wire   [3:1] MCInst_MC0_v0_3;
  wire   [3:0] MCInst_MC0_v0_2;
  wire   [3:1] MCInst_MC0_v0_1;
  wire   [2:1] MCInst_MC0_v0_0;
  wire   [3:0] MCInst_MC1_v3_3;
  wire   [3:0] MCInst_MC1_v3_2;
  wire   [3:0] MCInst_MC1_v3_1;
  wire   [3:1] MCInst_MC1_v3_0;
  wire   [3:0] MCInst_MC1_v2_3;
  wire   [3:0] MCInst_MC1_v2_2;
  wire   [3:0] MCInst_MC1_v2_1;
  wire   [3:1] MCInst_MC1_v2_0;
  wire   [3:1] MCInst_MC1_v1_3;
  wire   [3:0] MCInst_MC1_v1_2;
  wire   [3:0] MCInst_MC1_v1_1;
  wire   [3:1] MCInst_MC1_v0_3;
  wire   [3:0] MCInst_MC1_v0_2;
  wire   [3:1] MCInst_MC1_v0_1;
  wire   [2:1] MCInst_MC1_v0_0;
  wire   [3:0] MCInst_MC2_v3_3;
  wire   [3:0] MCInst_MC2_v3_2;
  wire   [3:0] MCInst_MC2_v3_1;
  wire   [3:1] MCInst_MC2_v3_0;
  wire   [3:0] MCInst_MC2_v2_3;
  wire   [3:0] MCInst_MC2_v2_2;
  wire   [3:0] MCInst_MC2_v2_1;
  wire   [3:1] MCInst_MC2_v2_0;
  wire   [3:1] MCInst_MC2_v1_3;
  wire   [3:0] MCInst_MC2_v1_2;
  wire   [3:0] MCInst_MC2_v1_1;
  wire   [3:1] MCInst_MC2_v0_3;
  wire   [3:0] MCInst_MC2_v0_2;
  wire   [3:1] MCInst_MC2_v0_1;
  wire   [2:1] MCInst_MC2_v0_0;
  wire   [3:0] MCInst_MC3_v3_3;
  wire   [3:0] MCInst_MC3_v3_2;
  wire   [3:0] MCInst_MC3_v3_1;
  wire   [3:1] MCInst_MC3_v3_0;
  wire   [3:0] MCInst_MC3_v2_3;
  wire   [3:0] MCInst_MC3_v2_2;
  wire   [3:0] MCInst_MC3_v2_1;
  wire   [3:1] MCInst_MC3_v2_0;
  wire   [3:1] MCInst_MC3_v1_3;
  wire   [3:0] MCInst_MC3_v1_2;
  wire   [3:0] MCInst_MC3_v1_1;
  wire   [3:1] MCInst_MC3_v0_3;
  wire   [3:0] MCInst_MC3_v0_2;
  wire   [3:1] MCInst_MC3_v0_1;
  wire   [2:1] MCInst_MC3_v0_0;
  wire   [3:0] MCInst2_MC0_v3_3;
  wire   [3:0] MCInst2_MC0_v3_2;
  wire   [3:0] MCInst2_MC0_v3_1;
  wire   [3:1] MCInst2_MC0_v3_0;
  wire   [3:0] MCInst2_MC0_v2_3;
  wire   [3:0] MCInst2_MC0_v2_2;
  wire   [3:0] MCInst2_MC0_v2_1;
  wire   [3:1] MCInst2_MC0_v2_0;
  wire   [3:1] MCInst2_MC0_v1_3;
  wire   [3:0] MCInst2_MC0_v1_2;
  wire   [3:0] MCInst2_MC0_v1_1;
  wire   [3:1] MCInst2_MC0_v0_3;
  wire   [3:0] MCInst2_MC0_v0_2;
  wire   [3:1] MCInst2_MC0_v0_1;
  wire   [2:1] MCInst2_MC0_v0_0;
  wire   [3:0] MCInst2_MC1_v3_3;
  wire   [3:0] MCInst2_MC1_v3_2;
  wire   [3:0] MCInst2_MC1_v3_1;
  wire   [3:1] MCInst2_MC1_v3_0;
  wire   [3:0] MCInst2_MC1_v2_3;
  wire   [3:0] MCInst2_MC1_v2_2;
  wire   [3:0] MCInst2_MC1_v2_1;
  wire   [3:1] MCInst2_MC1_v2_0;
  wire   [3:1] MCInst2_MC1_v1_3;
  wire   [3:0] MCInst2_MC1_v1_2;
  wire   [3:0] MCInst2_MC1_v1_1;
  wire   [3:1] MCInst2_MC1_v0_3;
  wire   [3:0] MCInst2_MC1_v0_2;
  wire   [3:1] MCInst2_MC1_v0_1;
  wire   [2:1] MCInst2_MC1_v0_0;
  wire   [3:0] MCInst2_MC2_v3_3;
  wire   [3:0] MCInst2_MC2_v3_2;
  wire   [3:0] MCInst2_MC2_v3_1;
  wire   [3:1] MCInst2_MC2_v3_0;
  wire   [3:0] MCInst2_MC2_v2_3;
  wire   [3:0] MCInst2_MC2_v2_2;
  wire   [3:0] MCInst2_MC2_v2_1;
  wire   [3:1] MCInst2_MC2_v2_0;
  wire   [3:1] MCInst2_MC2_v1_3;
  wire   [3:0] MCInst2_MC2_v1_2;
  wire   [3:0] MCInst2_MC2_v1_1;
  wire   [3:1] MCInst2_MC2_v0_3;
  wire   [3:0] MCInst2_MC2_v0_2;
  wire   [3:1] MCInst2_MC2_v0_1;
  wire   [2:1] MCInst2_MC2_v0_0;
  wire   [3:0] MCInst2_MC3_v3_3;
  wire   [3:0] MCInst2_MC3_v3_2;
  wire   [3:0] MCInst2_MC3_v3_1;
  wire   [3:1] MCInst2_MC3_v3_0;
  wire   [3:0] MCInst2_MC3_v2_3;
  wire   [3:0] MCInst2_MC3_v2_2;
  wire   [3:0] MCInst2_MC3_v2_1;
  wire   [3:1] MCInst2_MC3_v2_0;
  wire   [3:1] MCInst2_MC3_v1_3;
  wire   [3:0] MCInst2_MC3_v1_2;
  wire   [3:0] MCInst2_MC3_v1_1;
  wire   [3:1] MCInst2_MC3_v0_3;
  wire   [3:0] MCInst2_MC3_v0_2;
  wire   [3:1] MCInst2_MC3_v0_1;
  wire   [2:1] MCInst2_MC3_v0_0;
  wire   [2:0] Red_MCInst_MC0_v3_3;
  wire   [2:0] Red_MCInst_MC0_v3_2;
  wire   [2:1] Red_MCInst_MC0_v3_1;
  wire   [2:0] Red_MCInst_MC0_v3_0;
  wire   [2:0] Red_MCInst_MC0_v2_3;
  wire   [2:0] Red_MCInst_MC0_v2_2;
  wire   [2:0] Red_MCInst_MC0_v2_1;
  wire   [2:0] Red_MCInst_MC0_v2_0;
  wire   [2:0] Red_MCInst_MC0_v1_3;
  wire   [2:0] Red_MCInst_MC0_v1_2;
  wire   [2:1] Red_MCInst_MC0_v1_1;
  wire   [2:0] Red_MCInst_MC0_v1_0;
  wire   [2:0] Red_MCInst_MC0_v0_3;
  wire   [2:0] Red_MCInst_MC0_v0_2;
  wire   [2:0] Red_MCInst_MC0_v0_1;
  wire   [2:0] Red_MCInst_MC0_v0_0;
  wire   [2:0] Red_MCInst_MC1_v3_3;
  wire   [2:0] Red_MCInst_MC1_v3_2;
  wire   [2:1] Red_MCInst_MC1_v3_1;
  wire   [2:0] Red_MCInst_MC1_v3_0;
  wire   [2:0] Red_MCInst_MC1_v2_3;
  wire   [2:0] Red_MCInst_MC1_v2_2;
  wire   [2:0] Red_MCInst_MC1_v2_1;
  wire   [2:0] Red_MCInst_MC1_v2_0;
  wire   [2:0] Red_MCInst_MC1_v1_3;
  wire   [2:0] Red_MCInst_MC1_v1_2;
  wire   [2:1] Red_MCInst_MC1_v1_1;
  wire   [2:0] Red_MCInst_MC1_v1_0;
  wire   [2:0] Red_MCInst_MC1_v0_3;
  wire   [2:0] Red_MCInst_MC1_v0_2;
  wire   [2:0] Red_MCInst_MC1_v0_1;
  wire   [2:0] Red_MCInst_MC1_v0_0;
  wire   [2:0] Red_MCInst_MC2_v3_3;
  wire   [2:0] Red_MCInst_MC2_v3_2;
  wire   [2:1] Red_MCInst_MC2_v3_1;
  wire   [2:0] Red_MCInst_MC2_v3_0;
  wire   [2:0] Red_MCInst_MC2_v2_3;
  wire   [2:0] Red_MCInst_MC2_v2_2;
  wire   [2:0] Red_MCInst_MC2_v2_1;
  wire   [2:0] Red_MCInst_MC2_v2_0;
  wire   [2:0] Red_MCInst_MC2_v1_3;
  wire   [2:0] Red_MCInst_MC2_v1_2;
  wire   [2:1] Red_MCInst_MC2_v1_1;
  wire   [2:0] Red_MCInst_MC2_v1_0;
  wire   [2:0] Red_MCInst_MC2_v0_3;
  wire   [2:0] Red_MCInst_MC2_v0_2;
  wire   [2:0] Red_MCInst_MC2_v0_1;
  wire   [2:0] Red_MCInst_MC2_v0_0;
  wire   [2:0] Red_MCInst_MC3_v3_3;
  wire   [2:0] Red_MCInst_MC3_v3_2;
  wire   [2:1] Red_MCInst_MC3_v3_1;
  wire   [2:0] Red_MCInst_MC3_v3_0;
  wire   [2:0] Red_MCInst_MC3_v2_3;
  wire   [2:0] Red_MCInst_MC3_v2_2;
  wire   [2:0] Red_MCInst_MC3_v2_1;
  wire   [2:0] Red_MCInst_MC3_v2_0;
  wire   [2:0] Red_MCInst_MC3_v1_3;
  wire   [2:0] Red_MCInst_MC3_v1_2;
  wire   [2:1] Red_MCInst_MC3_v1_1;
  wire   [2:0] Red_MCInst_MC3_v1_0;
  wire   [2:0] Red_MCInst_MC3_v0_3;
  wire   [2:0] Red_MCInst_MC3_v0_2;
  wire   [2:0] Red_MCInst_MC3_v0_1;
  wire   [2:0] Red_MCInst_MC3_v0_0;
  wire   [2:0] Red_MCInst2_MC0_v3_3;
  wire   [2:0] Red_MCInst2_MC0_v3_2;
  wire   [2:1] Red_MCInst2_MC0_v3_1;
  wire   [2:0] Red_MCInst2_MC0_v3_0;
  wire   [2:0] Red_MCInst2_MC0_v2_3;
  wire   [2:0] Red_MCInst2_MC0_v2_2;
  wire   [2:0] Red_MCInst2_MC0_v2_1;
  wire   [2:0] Red_MCInst2_MC0_v2_0;
  wire   [2:0] Red_MCInst2_MC0_v1_3;
  wire   [2:0] Red_MCInst2_MC0_v1_2;
  wire   [2:1] Red_MCInst2_MC0_v1_1;
  wire   [2:0] Red_MCInst2_MC0_v1_0;
  wire   [2:0] Red_MCInst2_MC0_v0_3;
  wire   [2:0] Red_MCInst2_MC0_v0_2;
  wire   [2:0] Red_MCInst2_MC0_v0_1;
  wire   [2:0] Red_MCInst2_MC0_v0_0;
  wire   [2:0] Red_MCInst2_MC1_v3_3;
  wire   [2:0] Red_MCInst2_MC1_v3_2;
  wire   [2:1] Red_MCInst2_MC1_v3_1;
  wire   [2:0] Red_MCInst2_MC1_v3_0;
  wire   [2:0] Red_MCInst2_MC1_v2_3;
  wire   [2:0] Red_MCInst2_MC1_v2_2;
  wire   [2:0] Red_MCInst2_MC1_v2_1;
  wire   [2:0] Red_MCInst2_MC1_v2_0;
  wire   [2:0] Red_MCInst2_MC1_v1_3;
  wire   [2:0] Red_MCInst2_MC1_v1_2;
  wire   [2:1] Red_MCInst2_MC1_v1_1;
  wire   [2:0] Red_MCInst2_MC1_v1_0;
  wire   [2:0] Red_MCInst2_MC1_v0_3;
  wire   [2:0] Red_MCInst2_MC1_v0_2;
  wire   [2:0] Red_MCInst2_MC1_v0_1;
  wire   [2:0] Red_MCInst2_MC1_v0_0;
  wire   [2:0] Red_MCInst2_MC2_v3_3;
  wire   [2:0] Red_MCInst2_MC2_v3_2;
  wire   [2:1] Red_MCInst2_MC2_v3_1;
  wire   [2:0] Red_MCInst2_MC2_v3_0;
  wire   [2:0] Red_MCInst2_MC2_v2_3;
  wire   [2:0] Red_MCInst2_MC2_v2_2;
  wire   [2:0] Red_MCInst2_MC2_v2_1;
  wire   [2:0] Red_MCInst2_MC2_v2_0;
  wire   [2:0] Red_MCInst2_MC2_v1_3;
  wire   [2:0] Red_MCInst2_MC2_v1_2;
  wire   [2:1] Red_MCInst2_MC2_v1_1;
  wire   [2:0] Red_MCInst2_MC2_v1_0;
  wire   [2:0] Red_MCInst2_MC2_v0_3;
  wire   [2:0] Red_MCInst2_MC2_v0_2;
  wire   [2:0] Red_MCInst2_MC2_v0_1;
  wire   [2:0] Red_MCInst2_MC2_v0_0;
  wire   [2:0] Red_MCInst2_MC3_v3_3;
  wire   [2:0] Red_MCInst2_MC3_v3_2;
  wire   [2:1] Red_MCInst2_MC3_v3_1;
  wire   [2:0] Red_MCInst2_MC3_v3_0;
  wire   [2:0] Red_MCInst2_MC3_v2_3;
  wire   [2:0] Red_MCInst2_MC3_v2_2;
  wire   [2:0] Red_MCInst2_MC3_v2_1;
  wire   [2:0] Red_MCInst2_MC3_v2_0;
  wire   [2:0] Red_MCInst2_MC3_v1_3;
  wire   [2:0] Red_MCInst2_MC3_v1_2;
  wire   [2:1] Red_MCInst2_MC3_v1_1;
  wire   [2:0] Red_MCInst2_MC3_v1_0;
  wire   [2:0] Red_MCInst2_MC3_v0_3;
  wire   [2:0] Red_MCInst2_MC3_v0_2;
  wire   [2:0] Red_MCInst2_MC3_v0_1;
  wire   [2:0] Red_MCInst2_MC3_v0_0;

  AND2_X1 U6 ( .A1(Error[1]), .A2(Error[2]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(Error[0]), .A2(n4), .ZN(ErrorFlag) );
  XOR2_X2 AddKeyXOR_XORInst_0_0_U1 ( .A(Plaintext[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X2 AddKeyXOR_XORInst_0_1_U1 ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X2 AddKeyXOR_XORInst_0_2_U1 ( .A(Plaintext[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X2 AddKeyXOR_XORInst_0_3_U1 ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X2 AddKeyXOR_XORInst_1_0_U1 ( .A(Plaintext[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X2 AddKeyXOR_XORInst_1_1_U1 ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X2 AddKeyXOR_XORInst_1_2_U1 ( .A(Plaintext[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X2 AddKeyXOR_XORInst_1_3_U1 ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X2 AddKeyXOR_XORInst_2_0_U1 ( .A(Plaintext[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X2 AddKeyXOR_XORInst_2_1_U1 ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X2 AddKeyXOR_XORInst_2_2_U1 ( .A(Plaintext[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X2 AddKeyXOR_XORInst_2_3_U1 ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X2 AddKeyXOR_XORInst_3_0_U1 ( .A(Plaintext[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X2 AddKeyXOR_XORInst_3_1_U1 ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X2 AddKeyXOR_XORInst_3_2_U1 ( .A(Plaintext[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X2 AddKeyXOR_XORInst_3_3_U1 ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X2 AddKeyXOR_XORInst_4_0_U1 ( .A(Plaintext[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X2 AddKeyXOR_XORInst_4_1_U1 ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X2 AddKeyXOR_XORInst_4_2_U1 ( .A(Plaintext[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X2 AddKeyXOR_XORInst_4_3_U1 ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X2 AddKeyXOR_XORInst_5_0_U1 ( .A(Plaintext[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X2 AddKeyXOR_XORInst_5_1_U1 ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X2 AddKeyXOR_XORInst_5_2_U1 ( .A(Plaintext[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X2 AddKeyXOR_XORInst_5_3_U1 ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X2 AddKeyXOR_XORInst_6_0_U1 ( .A(Plaintext[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X2 AddKeyXOR_XORInst_6_1_U1 ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X2 AddKeyXOR_XORInst_6_2_U1 ( .A(Plaintext[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X2 AddKeyXOR_XORInst_6_3_U1 ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X2 AddKeyXOR_XORInst_7_0_U1 ( .A(Plaintext[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X2 AddKeyXOR_XORInst_7_1_U1 ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X2 AddKeyXOR_XORInst_7_2_U1 ( .A(Plaintext[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X2 AddKeyXOR_XORInst_7_3_U1 ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X2 AddKeyXOR_XORInst_8_0_U1 ( .A(Plaintext[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X2 AddKeyXOR_XORInst_8_1_U1 ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X2 AddKeyXOR_XORInst_8_2_U1 ( .A(Plaintext[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X2 AddKeyXOR_XORInst_8_3_U1 ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X2 AddKeyXOR_XORInst_9_0_U1 ( .A(Plaintext[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X2 AddKeyXOR_XORInst_9_1_U1 ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X2 AddKeyXOR_XORInst_9_2_U1 ( .A(Plaintext[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X2 AddKeyXOR_XORInst_9_3_U1 ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  XOR2_X2 AddKeyXOR_XORInst_10_0_U1 ( .A(Plaintext[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X2 AddKeyXOR_XORInst_10_1_U1 ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X2 AddKeyXOR_XORInst_10_2_U1 ( .A(Plaintext[42]), .B(Key[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X2 AddKeyXOR_XORInst_10_3_U1 ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X2 AddKeyXOR_XORInst_11_0_U1 ( .A(Plaintext[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X2 AddKeyXOR_XORInst_11_1_U1 ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X2 AddKeyXOR_XORInst_11_2_U1 ( .A(Plaintext[46]), .B(Key[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X2 AddKeyXOR_XORInst_11_3_U1 ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X2 AddKeyXOR_XORInst_12_0_U1 ( .A(Plaintext[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X2 AddKeyXOR_XORInst_12_1_U1 ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X2 AddKeyXOR_XORInst_12_2_U1 ( .A(Plaintext[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X2 AddKeyXOR_XORInst_12_3_U1 ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X2 AddKeyXOR_XORInst_13_0_U1 ( .A(Plaintext[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X2 AddKeyXOR_XORInst_13_1_U1 ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X2 AddKeyXOR_XORInst_13_2_U1 ( .A(Plaintext[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X2 AddKeyXOR_XORInst_13_3_U1 ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X2 AddKeyXOR_XORInst_14_0_U1 ( .A(Plaintext[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X2 AddKeyXOR_XORInst_14_1_U1 ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X2 AddKeyXOR_XORInst_14_2_U1 ( .A(Plaintext[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X2 AddKeyXOR_XORInst_14_3_U1 ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X2 AddKeyXOR_XORInst_15_0_U1 ( .A(Plaintext[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X2 AddKeyXOR_XORInst_15_1_U1 ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X2 AddKeyXOR_XORInst_15_2_U1 ( .A(Plaintext[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X2 AddKeyXOR_XORInst_15_3_U1 ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_0_U5 ( .A1(AddRoundKeyOutput[2]), .A2(
        SubCellInst_LFInst_0_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U4 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U3 ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_0_LFInst_0_n10), .ZN(MCInst_MC0_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_0_LFInst_0_n9), .B(SubCellInst_LFInst_0_LFInst_0_n8), .Z(SubCellInst_LFInst_0_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n24), .A2(
        SubCellInst_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U9 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U8 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n21), .A2(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n20), .A2(
        SubCellInst_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U5 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n19), .A2(
        SubCellInst_LFInst_0_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U3 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U2 ( .A(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_0_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n26), .A2(
        SubCellInst_LFInst_0_LFInst_1_n25), .ZN(Red_MCInst_MC0_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n25), .A2(
        SubCellInst_LFInst_0_LFInst_2_n28), .ZN(MCInst_MC0_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U7 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_0_LFInst_2_n26), .B(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n22), .A2(
        SubCellInst_LFInst_0_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_2_U3 ( .A(AddRoundKeyOutput[2]), .B(
        SubCellInst_LFInst_0_LFInst_2_n23), .Z(
        SubCellInst_LFInst_0_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U9 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n23), .A2(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U7 ( .A1(AddRoundKeyOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n23), .A2(
        SubCellInst_LFInst_0_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n20), .A2(
        SubCellInst_LFInst_0_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4 ( .A1(AddRoundKeyOutput[2]), .A2(
        AddRoundKeyOutput[0]), .ZN(SubCellInst_LFInst_0_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_0_LFInst_3_U3 ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U2 ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n26), .A2(
        SubCellInst_LFInst_0_LFInst_3_n25), .ZN(Red_MCInst_MC0_v3_1[2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_0_U5 ( .A1(AddRoundKeyOutput[6]), .A2(
        SubCellInst_LFInst_1_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U4 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U3 ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_1_LFInst_0_n10), .ZN(MCInst_MC3_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_1_LFInst_0_n9), .B(SubCellInst_LFInst_1_LFInst_0_n8), .Z(SubCellInst_LFInst_1_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n24), .A2(
        SubCellInst_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U9 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U8 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n21), .A2(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n20), .A2(
        SubCellInst_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U5 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n19), .A2(
        SubCellInst_LFInst_1_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U3 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U2 ( .A(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_1_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n26), .A2(
        SubCellInst_LFInst_1_LFInst_1_n25), .ZN(Red_MCInst_MC3_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n25), .A2(
        SubCellInst_LFInst_1_LFInst_2_n28), .ZN(MCInst_MC3_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U7 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_1_LFInst_2_n26), .B(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n22), .A2(
        SubCellInst_LFInst_1_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_2_U3 ( .A(AddRoundKeyOutput[6]), .B(
        SubCellInst_LFInst_1_LFInst_2_n23), .Z(
        SubCellInst_LFInst_1_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U2 ( .A1(AddRoundKeyOutput[5]), .A2(
        AddRoundKeyOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U9 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n23), .A2(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U7 ( .A1(AddRoundKeyOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n23), .A2(
        SubCellInst_LFInst_1_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n20), .A2(
        SubCellInst_LFInst_1_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4 ( .A1(AddRoundKeyOutput[6]), .A2(
        AddRoundKeyOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_1_LFInst_3_U3 ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U2 ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n26), .A2(
        SubCellInst_LFInst_1_LFInst_3_n25), .ZN(Red_MCInst_MC3_v3_1[2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_0_U5 ( .A1(AddRoundKeyOutput[10]), .A2(
        SubCellInst_LFInst_2_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U4 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U3 ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .Z(SubCellInst_LFInst_2_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_2_LFInst_0_n10), .ZN(MCInst_MC2_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_2_LFInst_0_n9), .B(SubCellInst_LFInst_2_LFInst_0_n8), .Z(SubCellInst_LFInst_2_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n24), .A2(
        SubCellInst_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U9 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U8 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n21), .A2(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n20), .A2(
        SubCellInst_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U5 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n19), .A2(
        SubCellInst_LFInst_2_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U3 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U2 ( .A(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_2_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n26), .A2(
        SubCellInst_LFInst_2_LFInst_1_n25), .ZN(Red_MCInst_MC2_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n25), .A2(
        SubCellInst_LFInst_2_LFInst_2_n28), .ZN(MCInst_MC2_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U7 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_2_LFInst_2_n26), .B(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n22), .A2(
        SubCellInst_LFInst_2_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_2_U3 ( .A(AddRoundKeyOutput[10]), .B(
        SubCellInst_LFInst_2_LFInst_2_n23), .Z(
        SubCellInst_LFInst_2_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U2 ( .A1(AddRoundKeyOutput[9]), .A2(
        AddRoundKeyOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U1 ( .A(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U9 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n23), .A2(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U7 ( .A1(AddRoundKeyOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n23), .A2(
        SubCellInst_LFInst_2_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n20), .A2(
        SubCellInst_LFInst_2_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4 ( .A1(AddRoundKeyOutput[10]), .A2(
        AddRoundKeyOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_2_LFInst_3_U3 ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U2 ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n26), .A2(
        SubCellInst_LFInst_2_LFInst_3_n25), .ZN(Red_MCInst_MC2_v3_1[2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_0_U5 ( .A1(AddRoundKeyOutput[14]), .A2(
        SubCellInst_LFInst_3_LFInst_0_n7), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U4 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n7) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U3 ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .Z(SubCellInst_LFInst_3_LFInst_0_n9) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_3_LFInst_0_n10), .ZN(MCInst_MC1_v3_2[3]) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_3_LFInst_0_n9), .B(SubCellInst_LFInst_3_LFInst_0_n8), .Z(SubCellInst_LFInst_3_LFInst_0_n10) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n24), .A2(
        SubCellInst_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U9 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U8 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n21), .A2(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n20), .A2(
        SubCellInst_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U5 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n19), .A2(
        SubCellInst_LFInst_3_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U3 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U2 ( .A(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n19) );
  NAND2_X2 SubCellInst_LFInst_3_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n26), .A2(
        SubCellInst_LFInst_3_LFInst_1_n25), .ZN(Red_MCInst_MC1_v3_3[2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n25), .A2(
        SubCellInst_LFInst_3_LFInst_2_n28), .ZN(MCInst_MC1_v3_0[3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U7 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_3_LFInst_2_n26), .B(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n22), .A2(
        SubCellInst_LFInst_3_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_2_U3 ( .A(AddRoundKeyOutput[14]), .B(
        SubCellInst_LFInst_3_LFInst_2_n23), .Z(
        SubCellInst_LFInst_3_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U2 ( .A1(AddRoundKeyOutput[13]), .A2(
        AddRoundKeyOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U1 ( .A(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U9 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n23), .A2(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U7 ( .A1(AddRoundKeyOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n23), .A2(
        SubCellInst_LFInst_3_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n20), .A2(
        SubCellInst_LFInst_3_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4 ( .A1(AddRoundKeyOutput[14]), .A2(
        AddRoundKeyOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_3_LFInst_3_U3 ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U2 ( .A1(AddRoundKeyOutput[12]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n26), .A2(
        SubCellInst_LFInst_3_LFInst_3_n25), .ZN(Red_MCInst_MC1_v3_1[2]) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_4_LFInst_0_n8), .B(SubCellInst_LFInst_4_LFInst_0_n7), .ZN(ShiftRowsOutput[24]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(AddRoundKeyOutput[18]), .A2(
        SubCellInst_LFInst_4_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U2 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n24), .A2(
        SubCellInst_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U9 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U8 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n21), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n20), .A2(
        SubCellInst_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U5 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n19), .A2(
        SubCellInst_LFInst_4_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U3 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U2 ( .A(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n26), .A2(
        SubCellInst_LFInst_4_LFInst_1_n25), .ZN(MCInst_MC1_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U9 ( .A1(AddRoundKeyOutput[18]), .A2(
        SubCellInst_LFInst_4_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_2_U8 ( .A1(AddRoundKeyOutput[17]), .A2(
        SubCellInst_LFInst_4_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U7 ( .A(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n25), .A2(
        SubCellInst_LFInst_4_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_4_LFInst_2_n23), .B(AddRoundKeyOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n22), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_2_U2 ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_4_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n29), .A2(
        SubCellInst_LFInst_4_LFInst_2_n28), .ZN(MCInst_MC1_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n25), .A2(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n25), .A2(
        SubCellInst_LFInst_4_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n22), .A2(
        SubCellInst_LFInst_4_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U6 ( .A1(AddRoundKeyOutput[18]), .A2(
        AddRoundKeyOutput[16]), .ZN(SubCellInst_LFInst_4_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_4_LFInst_3_U5 ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4 ( .A1(AddRoundKeyOutput[16]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_3_U3 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U2 ( .A1(AddRoundKeyOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_4_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n19), .A2(
        SubCellInst_LFInst_4_LFInst_3_n20), .ZN(Red_MCInst_MC1_v2_2[1]) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_5_LFInst_0_n8), .B(SubCellInst_LFInst_5_LFInst_0_n7), .ZN(ShiftRowsOutput[28]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(AddRoundKeyOutput[22]), .A2(
        SubCellInst_LFInst_5_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U2 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n24), .A2(
        SubCellInst_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U9 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U8 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n21), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n20), .A2(
        SubCellInst_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U5 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n19), .A2(
        SubCellInst_LFInst_5_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U3 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U2 ( .A(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n26), .A2(
        SubCellInst_LFInst_5_LFInst_1_n25), .ZN(MCInst_MC0_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U9 ( .A1(AddRoundKeyOutput[22]), .A2(
        SubCellInst_LFInst_5_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_2_U8 ( .A1(AddRoundKeyOutput[21]), .A2(
        SubCellInst_LFInst_5_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U7 ( .A(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n25), .A2(
        SubCellInst_LFInst_5_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_5_LFInst_2_n23), .B(AddRoundKeyOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n22), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_2_U2 ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_5_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n29), .A2(
        SubCellInst_LFInst_5_LFInst_2_n28), .ZN(MCInst_MC0_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n25), .A2(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n25), .A2(
        SubCellInst_LFInst_5_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n22), .A2(
        SubCellInst_LFInst_5_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U6 ( .A1(AddRoundKeyOutput[22]), .A2(
        AddRoundKeyOutput[20]), .ZN(SubCellInst_LFInst_5_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_5_LFInst_3_U5 ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4 ( .A1(AddRoundKeyOutput[20]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_3_U3 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U2 ( .A1(AddRoundKeyOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_5_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n19), .A2(
        SubCellInst_LFInst_5_LFInst_3_n20), .ZN(Red_MCInst_MC0_v2_2[1]) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_6_LFInst_0_n8), .B(SubCellInst_LFInst_6_LFInst_0_n7), .ZN(ShiftRowsOutput[16]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(AddRoundKeyOutput[26]), .A2(
        SubCellInst_LFInst_6_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U2 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .Z(SubCellInst_LFInst_6_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n24), .A2(
        SubCellInst_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U9 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U8 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n21), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n20), .A2(
        SubCellInst_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U5 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n19), .A2(
        SubCellInst_LFInst_6_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U3 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U2 ( .A(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n26), .A2(
        SubCellInst_LFInst_6_LFInst_1_n25), .ZN(MCInst_MC3_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U9 ( .A1(AddRoundKeyOutput[26]), .A2(
        SubCellInst_LFInst_6_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_2_U8 ( .A1(AddRoundKeyOutput[25]), .A2(
        SubCellInst_LFInst_6_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U7 ( .A(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n25), .A2(
        SubCellInst_LFInst_6_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_6_LFInst_2_n23), .B(AddRoundKeyOutput[26]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n22), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_2_U2 ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_6_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n29), .A2(
        SubCellInst_LFInst_6_LFInst_2_n28), .ZN(MCInst_MC3_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n25), .A2(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n25), .A2(
        SubCellInst_LFInst_6_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n22), .A2(
        SubCellInst_LFInst_6_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U6 ( .A1(AddRoundKeyOutput[26]), .A2(
        AddRoundKeyOutput[24]), .ZN(SubCellInst_LFInst_6_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_6_LFInst_3_U5 ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4 ( .A1(AddRoundKeyOutput[24]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_3_U3 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U2 ( .A1(AddRoundKeyOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_6_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n19), .A2(
        SubCellInst_LFInst_6_LFInst_3_n20), .ZN(Red_MCInst_MC3_v2_2[1]) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_0_U4 ( .A(
        SubCellInst_LFInst_7_LFInst_0_n8), .B(SubCellInst_LFInst_7_LFInst_0_n7), .ZN(ShiftRowsOutput[20]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(AddRoundKeyOutput[30]), .A2(
        SubCellInst_LFInst_7_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U2 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .Z(SubCellInst_LFInst_7_LFInst_0_n8) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n24), .A2(
        SubCellInst_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U9 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U8 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n21), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n20), .A2(
        SubCellInst_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U5 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n19), .A2(
        SubCellInst_LFInst_7_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U3 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U2 ( .A(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n26), .A2(
        SubCellInst_LFInst_7_LFInst_1_n25), .ZN(MCInst_MC2_v2_0[2]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U9 ( .A1(AddRoundKeyOutput[30]), .A2(
        SubCellInst_LFInst_7_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n28) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_2_U8 ( .A1(AddRoundKeyOutput[29]), .A2(
        SubCellInst_LFInst_7_LFInst_2_n26), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n27) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U7 ( .A(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n25), .A2(
        SubCellInst_LFInst_7_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n29) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_2_U5 ( .A(
        SubCellInst_LFInst_7_LFInst_2_n23), .B(AddRoundKeyOutput[30]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n23) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n22), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n25) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_2_U2 ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n22) );
  NAND2_X2 SubCellInst_LFInst_7_LFInst_2_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n29), .A2(
        SubCellInst_LFInst_7_LFInst_2_n28), .ZN(MCInst_MC2_v2_0[3]) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U9 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n25), .A2(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n25), .A2(
        SubCellInst_LFInst_7_LFInst_3_n23), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n24) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U7 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n22), .A2(
        SubCellInst_LFInst_7_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n23) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U6 ( .A1(AddRoundKeyOutput[30]), .A2(
        AddRoundKeyOutput[28]), .ZN(SubCellInst_LFInst_7_LFInst_3_n21) );
  INV_X1 SubCellInst_LFInst_7_LFInst_3_U5 ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4 ( .A1(AddRoundKeyOutput[28]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_3_n25) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_3_U3 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n26), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U2 ( .A1(AddRoundKeyOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n19) );
  OR2_X2 SubCellInst_LFInst_7_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n19), .A2(
        SubCellInst_LFInst_7_LFInst_3_n20), .ZN(Red_MCInst_MC2_v2_2[1]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_0_U5 ( .A1(AddRoundKeyOutput[34]), .A2(
        SubCellInst_LFInst_8_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U4 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U3 ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_8_LFInst_0_n12), .ZN(MCInst_MC2_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_8_LFInst_0_n11), .B(
        SubCellInst_LFInst_8_LFInst_0_n10), .Z(
        SubCellInst_LFInst_8_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n24), .A2(
        SubCellInst_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U9 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U8 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n21), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n20), .A2(
        SubCellInst_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U5 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n19), .A2(
        SubCellInst_LFInst_8_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U3 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U2 ( .A(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n26), .A2(
        SubCellInst_LFInst_8_LFInst_1_n25), .ZN(MCInst_MC2_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n25), .A2(
        SubCellInst_LFInst_8_LFInst_2_n28), .ZN(MCInst_MC2_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U7 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_8_LFInst_2_n26), .B(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_2_U5 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n22), .A2(
        SubCellInst_LFInst_8_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U3 ( .A(AddRoundKeyOutput[34]), .B(
        SubCellInst_LFInst_8_LFInst_2_n23), .Z(
        SubCellInst_LFInst_8_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U2 ( .A1(AddRoundKeyOutput[33]), .A2(
        AddRoundKeyOutput[32]), .ZN(SubCellInst_LFInst_8_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U1 ( .A(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U9 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n23), .A2(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U7 ( .A1(AddRoundKeyOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n23), .A2(
        SubCellInst_LFInst_8_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n20), .A2(
        SubCellInst_LFInst_8_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U4 ( .A1(AddRoundKeyOutput[34]), .A2(
        AddRoundKeyOutput[32]), .ZN(SubCellInst_LFInst_8_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_8_LFInst_3_U3 ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U2 ( .A1(AddRoundKeyOutput[32]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n26), .A2(
        SubCellInst_LFInst_8_LFInst_3_n25), .ZN(Red_MCInst_MC2_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_0_U5 ( .A1(AddRoundKeyOutput[38]), .A2(
        SubCellInst_LFInst_9_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U4 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U3 ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_9_LFInst_0_n12), .ZN(MCInst_MC1_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_9_LFInst_0_n11), .B(
        SubCellInst_LFInst_9_LFInst_0_n10), .Z(
        SubCellInst_LFInst_9_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n24), .A2(
        SubCellInst_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U9 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U8 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n21), .A2(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n20), .A2(
        SubCellInst_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U5 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n19), .A2(
        SubCellInst_LFInst_9_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U3 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U2 ( .A(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n26), .A2(
        SubCellInst_LFInst_9_LFInst_1_n25), .ZN(MCInst_MC1_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n25), .A2(
        SubCellInst_LFInst_9_LFInst_2_n28), .ZN(MCInst_MC1_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U7 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_9_LFInst_2_n26), .B(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n22), .A2(
        SubCellInst_LFInst_9_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_2_U3 ( .A(AddRoundKeyOutput[38]), .B(
        SubCellInst_LFInst_9_LFInst_2_n23), .Z(
        SubCellInst_LFInst_9_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U2 ( .A1(AddRoundKeyOutput[37]), .A2(
        AddRoundKeyOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U1 ( .A(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U9 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n23), .A2(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U7 ( .A1(AddRoundKeyOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n23), .A2(
        SubCellInst_LFInst_9_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n20), .A2(
        SubCellInst_LFInst_9_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U4 ( .A1(AddRoundKeyOutput[38]), .A2(
        AddRoundKeyOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_9_LFInst_3_U3 ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U2 ( .A1(AddRoundKeyOutput[36]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n26), .A2(
        SubCellInst_LFInst_9_LFInst_3_n25), .ZN(Red_MCInst_MC1_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_0_U5 ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U4 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U3 ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .Z(SubCellInst_LFInst_10_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_10_LFInst_0_n12), .ZN(MCInst_MC0_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_10_LFInst_0_n11), .B(
        SubCellInst_LFInst_10_LFInst_0_n10), .Z(
        SubCellInst_LFInst_10_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n24), .A2(
        SubCellInst_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U9 ( .A1(AddRoundKeyOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U8 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n21), .A2(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n20), .A2(
        SubCellInst_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U5 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n19), .A2(
        SubCellInst_LFInst_10_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U3 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U2 ( .A(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n26), .A2(
        SubCellInst_LFInst_10_LFInst_1_n25), .ZN(MCInst_MC0_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n25), .A2(
        SubCellInst_LFInst_10_LFInst_2_n28), .ZN(MCInst_MC0_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U7 ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_10_LFInst_2_n26), .B(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(AddRoundKeyOutput[40]), .A2(
        AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n22), .A2(
        SubCellInst_LFInst_10_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_2_U3 ( .A(AddRoundKeyOutput[42]), .B(
        SubCellInst_LFInst_10_LFInst_2_n23), .Z(
        SubCellInst_LFInst_10_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U2 ( .A1(AddRoundKeyOutput[41]), 
        .A2(AddRoundKeyOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U1 ( .A(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U9 ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n23), .A2(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U7 ( .A1(AddRoundKeyOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n23), .A2(
        SubCellInst_LFInst_10_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n20), .A2(
        SubCellInst_LFInst_10_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U4 ( .A1(AddRoundKeyOutput[42]), .A2(
        AddRoundKeyOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_10_LFInst_3_U3 ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U2 ( .A1(AddRoundKeyOutput[40]), .A2(
        AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n26), .A2(
        SubCellInst_LFInst_10_LFInst_3_n25), .ZN(Red_MCInst_MC0_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_0_U5 ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_0_n9), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n10) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U4 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n9) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U3 ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .Z(SubCellInst_LFInst_11_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_11_LFInst_0_n12), .ZN(MCInst_MC3_v1_0_0_) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_11_LFInst_0_n11), .B(
        SubCellInst_LFInst_11_LFInst_0_n10), .Z(
        SubCellInst_LFInst_11_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n24), .A2(
        SubCellInst_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U9 ( .A1(AddRoundKeyOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U8 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n21), .A2(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n20), .A2(
        SubCellInst_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U5 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n19), .A2(
        SubCellInst_LFInst_11_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U3 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U2 ( .A(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n26), .A2(
        SubCellInst_LFInst_11_LFInst_1_n25), .ZN(MCInst_MC3_v1_3[2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n25), .A2(
        SubCellInst_LFInst_11_LFInst_2_n28), .ZN(MCInst_MC3_v1_3[3]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U7 ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_11_LFInst_2_n26), .B(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(AddRoundKeyOutput[44]), .A2(
        AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n22), .A2(
        SubCellInst_LFInst_11_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_2_U3 ( .A(AddRoundKeyOutput[46]), .B(
        SubCellInst_LFInst_11_LFInst_2_n23), .Z(
        SubCellInst_LFInst_11_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U2 ( .A1(AddRoundKeyOutput[45]), 
        .A2(AddRoundKeyOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U9 ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n23), .A2(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U7 ( .A1(AddRoundKeyOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n23), .A2(
        SubCellInst_LFInst_11_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n20), .A2(
        SubCellInst_LFInst_11_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U4 ( .A1(AddRoundKeyOutput[46]), .A2(
        AddRoundKeyOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_11_LFInst_3_U3 ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U2 ( .A1(AddRoundKeyOutput[44]), .A2(
        AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n26), .A2(
        SubCellInst_LFInst_11_LFInst_3_n25), .ZN(Red_MCInst_MC3_v1_1[2]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_0_U5 ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U4 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U3 ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_12_LFInst_0_n9), .ZN(Red_MCInst_MC3_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_12_LFInst_0_n8), .B(
        SubCellInst_LFInst_12_LFInst_0_n7), .Z(
        SubCellInst_LFInst_12_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n24), .A2(
        SubCellInst_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U9 ( .A1(AddRoundKeyOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U8 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n21), .A2(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n20), .A2(
        SubCellInst_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U5 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n19), .A2(
        SubCellInst_LFInst_12_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U3 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U2 ( .A(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n26), .A2(
        SubCellInst_LFInst_12_LFInst_1_n25), .ZN(Red_MCInst_MC3_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n25), .A2(
        SubCellInst_LFInst_12_LFInst_2_n28), .ZN(MCInst_MC3_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U7 ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_12_LFInst_2_n26), .B(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_2_U5 ( .A1(AddRoundKeyOutput[48]), .A2(
        AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n22), .A2(
        SubCellInst_LFInst_12_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U3 ( .A(AddRoundKeyOutput[50]), .B(
        SubCellInst_LFInst_12_LFInst_2_n23), .Z(
        SubCellInst_LFInst_12_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U2 ( .A1(AddRoundKeyOutput[49]), 
        .A2(AddRoundKeyOutput[48]), .ZN(SubCellInst_LFInst_12_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U1 ( .A(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U9 ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n23), .A2(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U7 ( .A1(AddRoundKeyOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n23), .A2(
        SubCellInst_LFInst_12_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n20), .A2(
        SubCellInst_LFInst_12_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U4 ( .A1(AddRoundKeyOutput[50]), .A2(
        AddRoundKeyOutput[48]), .ZN(SubCellInst_LFInst_12_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_12_LFInst_3_U3 ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U2 ( .A1(AddRoundKeyOutput[48]), .A2(
        AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n26), .A2(
        SubCellInst_LFInst_12_LFInst_3_n25), .ZN(Red_MCInst_MC3_v0_1[0]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_0_U5 ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U4 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U3 ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_13_LFInst_0_n9), .ZN(Red_MCInst_MC2_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_13_LFInst_0_n8), .B(
        SubCellInst_LFInst_13_LFInst_0_n7), .Z(
        SubCellInst_LFInst_13_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n24), .A2(
        SubCellInst_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U9 ( .A1(AddRoundKeyOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U8 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n21), .A2(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n20), .A2(
        SubCellInst_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U5 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n19), .A2(
        SubCellInst_LFInst_13_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U2 ( .A(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n26), .A2(
        SubCellInst_LFInst_13_LFInst_1_n25), .ZN(Red_MCInst_MC2_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n25), .A2(
        SubCellInst_LFInst_13_LFInst_2_n28), .ZN(MCInst_MC2_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U7 ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_13_LFInst_2_n26), .B(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_2_U5 ( .A1(AddRoundKeyOutput[52]), .A2(
        AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n22), .A2(
        SubCellInst_LFInst_13_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_2_U3 ( .A(AddRoundKeyOutput[54]), .B(
        SubCellInst_LFInst_13_LFInst_2_n23), .Z(
        SubCellInst_LFInst_13_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U2 ( .A1(AddRoundKeyOutput[53]), 
        .A2(AddRoundKeyOutput[52]), .ZN(SubCellInst_LFInst_13_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U9 ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n23), .A2(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U7 ( .A1(AddRoundKeyOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n23), .A2(
        SubCellInst_LFInst_13_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n20), .A2(
        SubCellInst_LFInst_13_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U4 ( .A1(AddRoundKeyOutput[54]), .A2(
        AddRoundKeyOutput[52]), .ZN(SubCellInst_LFInst_13_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_13_LFInst_3_U3 ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U2 ( .A1(AddRoundKeyOutput[52]), .A2(
        AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n26), .A2(
        SubCellInst_LFInst_13_LFInst_3_n25), .ZN(Red_MCInst_MC2_v0_1[0]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_0_U5 ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U4 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U3 ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .Z(SubCellInst_LFInst_14_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_14_LFInst_0_n9), .ZN(Red_MCInst_MC1_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_14_LFInst_0_n8), .B(
        SubCellInst_LFInst_14_LFInst_0_n7), .Z(
        SubCellInst_LFInst_14_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n24), .A2(
        SubCellInst_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U9 ( .A1(AddRoundKeyOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U8 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n21), .A2(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n20), .A2(
        SubCellInst_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U5 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n19), .A2(
        SubCellInst_LFInst_14_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U3 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U2 ( .A(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n26), .A2(
        SubCellInst_LFInst_14_LFInst_1_n25), .ZN(Red_MCInst_MC1_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n25), .A2(
        SubCellInst_LFInst_14_LFInst_2_n28), .ZN(MCInst_MC1_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U7 ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_14_LFInst_2_n26), .B(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_2_U5 ( .A1(AddRoundKeyOutput[56]), .A2(
        AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n22), .A2(
        SubCellInst_LFInst_14_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U3 ( .A(AddRoundKeyOutput[58]), .B(
        SubCellInst_LFInst_14_LFInst_2_n23), .Z(
        SubCellInst_LFInst_14_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U2 ( .A1(AddRoundKeyOutput[57]), 
        .A2(AddRoundKeyOutput[56]), .ZN(SubCellInst_LFInst_14_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U1 ( .A(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U9 ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n23), .A2(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U7 ( .A1(AddRoundKeyOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n23), .A2(
        SubCellInst_LFInst_14_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n20), .A2(
        SubCellInst_LFInst_14_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U4 ( .A1(AddRoundKeyOutput[58]), .A2(
        AddRoundKeyOutput[56]), .ZN(SubCellInst_LFInst_14_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_14_LFInst_3_U3 ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U2 ( .A1(AddRoundKeyOutput[56]), .A2(
        AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n26), .A2(
        SubCellInst_LFInst_14_LFInst_3_n25), .ZN(Red_MCInst_MC1_v0_1[0]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_0_U5 ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_0_n6), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n7) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U4 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n6) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U3 ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .Z(SubCellInst_LFInst_15_LFInst_0_n8) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U2 ( .A(
        SubCellInst_LFInst_15_LFInst_0_n9), .ZN(Red_MCInst_MC0_v0_0[0]) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U1 ( .A(
        SubCellInst_LFInst_15_LFInst_0_n8), .B(
        SubCellInst_LFInst_15_LFInst_0_n7), .Z(
        SubCellInst_LFInst_15_LFInst_0_n9) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U10 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n24), .A2(
        SubCellInst_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n25) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U9 ( .A1(AddRoundKeyOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_1_n22), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n24) );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U8 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n22) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U7 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n21), .A2(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n26) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n20), .A2(
        SubCellInst_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n21) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U5 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n23) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n19), .A2(
        SubCellInst_LFInst_15_LFInst_1_n18), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n20) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U3 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_1_n18) );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U2 ( .A(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n19) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U1 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n26), .A2(
        SubCellInst_LFInst_15_LFInst_1_n25), .ZN(Red_MCInst_MC0_v0_2[2]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U8 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n25), .A2(
        SubCellInst_LFInst_15_LFInst_2_n28), .ZN(MCInst_MC0_v0_3[3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U7 ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n27), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n28) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_2_U6 ( .A(
        SubCellInst_LFInst_15_LFInst_2_n26), .B(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n27) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_2_U5 ( .A1(AddRoundKeyOutput[60]), .A2(
        AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_2_n26) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n22), .A2(
        SubCellInst_LFInst_15_LFInst_2_n24), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n25) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U3 ( .A(AddRoundKeyOutput[62]), .B(
        SubCellInst_LFInst_15_LFInst_2_n23), .Z(
        SubCellInst_LFInst_15_LFInst_2_n24) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U2 ( .A1(AddRoundKeyOutput[61]), 
        .A2(AddRoundKeyOutput[60]), .ZN(SubCellInst_LFInst_15_LFInst_2_n23) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U1 ( .A(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n22) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U9 ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_3_n24), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n25) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U8 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n23), .A2(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n24) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U7 ( .A1(AddRoundKeyOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_3_n22), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n26) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n23), .A2(
        SubCellInst_LFInst_15_LFInst_3_n21), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n22) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U5 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n20), .A2(
        SubCellInst_LFInst_15_LFInst_3_n19), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n21) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U4 ( .A1(AddRoundKeyOutput[62]), .A2(
        AddRoundKeyOutput[60]), .ZN(SubCellInst_LFInst_15_LFInst_3_n19) );
  INV_X1 SubCellInst_LFInst_15_LFInst_3_U3 ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n20) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U2 ( .A1(AddRoundKeyOutput[60]), .A2(
        AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_3_n23) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n26), .A2(
        SubCellInst_LFInst_15_LFInst_3_n25), .ZN(Red_MCInst_MC0_v0_1[0]) );
  BUF_X1 MCInst_MC0_U2 ( .A(ShiftRowsOutput[28]), .Z(MCInst_MC0_v2_3[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U2 ( .A(MCInst_MC0_v0_2Inst_0_n3), .B(
        Red_MCInst_MC0_v0_1[0]), .ZN(MCInst_MC0_v0_2[0]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .ZN(MCInst_MC0_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v1_1Inst_0_U1 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .Z(MCInst_MC0_v1_1[0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U2 ( .A(MCInst_MC0_v1_2Inst_0_n3), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_v1_2[0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v2_1Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(MCInst_MC0_v2_1[0]) );
  XOR2_X1 MCInst_MC0_v2_2Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(MCInst_MC0_v2_2[0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U3 ( .A(MCInst_MC0_v2_3Inst_0_n6), .B(
        MCInst_MC0_v2_3Inst_0_n5), .ZN(MCInst_MC0_v2_3[0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC0_v2_3Inst_0_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC0_v3_1Inst_0_U1 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_v3_1[0]) );
  XOR2_X1 MCInst_MC0_v3_2Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_v3_2[0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U2 ( .A(MCInst_MC0_v3_3Inst_0_n3), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(MCInst_MC0_v3_3[0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(MCInst_MC0_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC0_v0_0Inst_1_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_0[1]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_1_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v0_3[3]), .Z(MCInst_MC0_v0_1[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U2 ( .A(MCInst_MC0_v0_2Inst_1_n3), .B(
        Red_MCInst_MC0_v0_1[0]), .ZN(MCInst_MC0_v0_2[1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .ZN(MCInst_MC0_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_3[1]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[3]), .Z(MCInst_MC0_v1_1[1]) );
  XOR2_X1 MCInst_MC0_v1_2Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .Z(MCInst_MC0_v1_2[1]) );
  XOR2_X1 MCInst_MC0_v1_3Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_1[2]), .Z(MCInst_MC0_v1_3[1]) );
  XOR2_X1 MCInst_MC0_v2_0Inst_1_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(MCInst_MC0_v2_0[1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U2 ( .A(MCInst_MC0_v2_1Inst_1_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_1[1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U3 ( .A(MCInst_MC0_v2_2Inst_1_n6), .B(
        MCInst_MC0_v2_2Inst_1_n5), .ZN(MCInst_MC0_v2_2[1]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC0_v2_2Inst_1_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC0_v3_0Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_v3_0[1]) );
  XOR2_X1 MCInst_MC0_v3_1Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_v3_1[1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U2 ( .A(MCInst_MC0_v3_3Inst_1_n3), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(MCInst_MC0_v3_3[1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .ZN(MCInst_MC0_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_0[2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_2_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_1[2]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_2[2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U2 ( .A(MCInst_MC0_v1_1Inst_2_n3), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_v1_1[2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U2 ( .A(MCInst_MC0_v1_2Inst_2_n3), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_v1_2[2]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U2 ( .A(MCInst_MC0_v2_1Inst_2_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_1[2]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U2 ( .A(MCInst_MC0_v2_2Inst_2_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_2[2]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC0_v2_3Inst_2_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(MCInst_MC0_v2_3[2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U2 ( .A(MCInst_MC0_v3_1Inst_2_n3), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(MCInst_MC0_v3_1[2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(MCInst_MC0_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC0_v3_3Inst_2_U1 ( .A(Red_MCInst_MC0_v3_3[2]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_v3_3[2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_3_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(MCInst_MC0_v0_1[3]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_3_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .Z(MCInst_MC0_v0_2[3]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_3_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        MCInst_MC0_v1_3[3]), .Z(MCInst_MC0_v1_1[3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U3 ( .A(MCInst_MC0_v1_2Inst_3_n6), .B(
        MCInst_MC0_v1_2Inst_3_n5), .ZN(MCInst_MC0_v1_2[3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U2 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC0_v1_2Inst_3_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .Z(MCInst_MC0_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC0_v2_1Inst_3_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(MCInst_MC0_v2_1[3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U2 ( .A(MCInst_MC0_v2_2Inst_3_n3), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(MCInst_MC0_v2_2[3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U2 ( .A(MCInst_MC0_v2_3Inst_3_n3), .B(
        MCInst_MC0_v2_0[3]), .ZN(MCInst_MC0_v2_3[3]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U1 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v2_0[2]), .ZN(MCInst_MC0_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC0_v3_1Inst_3_U1 ( .A(Red_MCInst_MC0_v3_3[2]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_v3_1[3]) );
  XOR2_X1 MCInst_MC0_v3_3Inst_3_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_v3_3[3]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_0_n8), .B(MCInst_MC0_r0Inst_XORInst_0_0_n7), .ZN(MC_output[60]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_2[1]), .B(
        MCInst_MC0_v1_0_0_), .ZN(MCInst_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_1_n8), .B(MCInst_MC0_r0Inst_XORInst_0_1_n7), .ZN(MC_output[61]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_0[1]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_0[1]), .B(
        MCInst_MC0_v3_0[1]), .Z(MCInst_MC0_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_2_n8), .B(MCInst_MC0_r0Inst_XORInst_0_2_n7), .ZN(MC_output[62]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_0[2]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r0Inst_XORInst_0_3_n8), .B(MCInst_MC0_r0Inst_XORInst_0_3_n7), .ZN(MC_output[63]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_0_n8), .B(MCInst_MC0_r1Inst_XORInst_0_0_n7), .ZN(MC_output[44]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_1[0]), .B(
        MCInst_MC0_v1_1[0]), .ZN(MCInst_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_1[0]), .Z(MCInst_MC0_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_1_n8), .B(MCInst_MC0_r1Inst_XORInst_0_1_n7), .ZN(MC_output[45]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v1_1[1]), .ZN(MCInst_MC0_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_1[1]), .B(
        MCInst_MC0_v3_1[1]), .Z(MCInst_MC0_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_2_n8), .B(MCInst_MC0_r1Inst_XORInst_0_2_n7), .ZN(MC_output[46]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_1[2]), .B(
        MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_1[2]), .B(
        MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r1Inst_XORInst_0_3_n8), .B(MCInst_MC0_r1Inst_XORInst_0_3_n7), .ZN(MC_output[47]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_1[3]), .B(
        MCInst_MC0_v1_1[3]), .ZN(MCInst_MC0_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_1[3]), .B(
        MCInst_MC0_v3_1[3]), .Z(MCInst_MC0_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_0_n8), .B(MCInst_MC0_r2Inst_XORInst_0_0_n7), .ZN(MC_output[28]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_2[0]), .B(
        MCInst_MC0_v1_2[0]), .ZN(MCInst_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC0_v0_2[0]), .B(
        MCInst_MC0_v3_2[0]), .Z(MCInst_MC0_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_1_n8), .B(MCInst_MC0_r2Inst_XORInst_0_1_n7), .ZN(MC_output[29]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_2[1]), .B(
        MCInst_MC0_v1_2[1]), .ZN(MCInst_MC0_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_2[1]), .B(
        MCInst_MC0_v3_0[3]), .Z(MCInst_MC0_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_2_n8), .B(MCInst_MC0_r2Inst_XORInst_0_2_n7), .ZN(MC_output[30]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_2[2]), .B(
        MCInst_MC0_v1_2[2]), .ZN(MCInst_MC0_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC0_v0_2[2]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(MCInst_MC0_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r2Inst_XORInst_0_3_n8), .B(MCInst_MC0_r2Inst_XORInst_0_3_n7), .ZN(MC_output[31]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_2[3]), .B(
        MCInst_MC0_v1_2[3]), .ZN(MCInst_MC0_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_2[3]), .B(
        MCInst_MC0_v3_2[3]), .Z(MCInst_MC0_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_0_n8), .B(MCInst_MC0_r3Inst_XORInst_0_0_n7), .ZN(MC_output[12]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC0_v2_3[0]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(MCInst_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_1[0]), .B(
        MCInst_MC0_v3_3[0]), .Z(MCInst_MC0_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_1_n8), .B(MCInst_MC0_r3Inst_XORInst_0_1_n7), .ZN(MC_output[13]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC0_v2_3[1]), .B(
        MCInst_MC0_v1_3[1]), .ZN(MCInst_MC0_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC0_v0_3[1]), .B(
        MCInst_MC0_v3_3[1]), .Z(MCInst_MC0_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_2_n8), .B(MCInst_MC0_r3Inst_XORInst_0_2_n7), .ZN(MC_output[14]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC0_v2_3[2]), .B(
        MCInst_MC0_v1_3[2]), .ZN(MCInst_MC0_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        MCInst_MC0_v3_3[2]), .Z(MCInst_MC0_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC0_r3Inst_XORInst_0_3_n8), .B(MCInst_MC0_r3Inst_XORInst_0_3_n7), .ZN(MC_output[15]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC0_v2_3[3]), .B(
        MCInst_MC0_v1_3[3]), .ZN(MCInst_MC0_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        MCInst_MC0_v3_3[3]), .Z(MCInst_MC0_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst_MC1_U2 ( .A(ShiftRowsOutput[24]), .Z(MCInst_MC1_v2_3[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U2 ( .A(MCInst_MC1_v0_2Inst_0_n3), .B(
        Red_MCInst_MC1_v0_1[0]), .ZN(MCInst_MC1_v0_2[0]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .ZN(MCInst_MC1_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v1_1Inst_0_U1 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .Z(MCInst_MC1_v1_1[0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U2 ( .A(MCInst_MC1_v1_2Inst_0_n3), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_v1_2[0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v2_1Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(MCInst_MC1_v2_1[0]) );
  XOR2_X1 MCInst_MC1_v2_2Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(MCInst_MC1_v2_2[0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U3 ( .A(MCInst_MC1_v2_3Inst_0_n6), .B(
        MCInst_MC1_v2_3Inst_0_n5), .ZN(MCInst_MC1_v2_3[0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC1_v2_3Inst_0_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC1_v3_1Inst_0_U1 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_v3_1[0]) );
  XOR2_X1 MCInst_MC1_v3_2Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_v3_2[0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U2 ( .A(MCInst_MC1_v3_3Inst_0_n3), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(MCInst_MC1_v3_3[0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(MCInst_MC1_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC1_v0_0Inst_1_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_0[1]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_1_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v0_3[3]), .Z(MCInst_MC1_v0_1[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U2 ( .A(MCInst_MC1_v0_2Inst_1_n3), .B(
        Red_MCInst_MC1_v0_1[0]), .ZN(MCInst_MC1_v0_2[1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .ZN(MCInst_MC1_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_3[1]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[3]), .Z(MCInst_MC1_v1_1[1]) );
  XOR2_X1 MCInst_MC1_v1_2Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .Z(MCInst_MC1_v1_2[1]) );
  XOR2_X1 MCInst_MC1_v1_3Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_1[2]), .Z(MCInst_MC1_v1_3[1]) );
  XOR2_X1 MCInst_MC1_v2_0Inst_1_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(MCInst_MC1_v2_0[1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U2 ( .A(MCInst_MC1_v2_1Inst_1_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_1[1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U3 ( .A(MCInst_MC1_v2_2Inst_1_n6), .B(
        MCInst_MC1_v2_2Inst_1_n5), .ZN(MCInst_MC1_v2_2[1]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC1_v2_2Inst_1_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC1_v3_0Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_v3_0[1]) );
  XOR2_X1 MCInst_MC1_v3_1Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_v3_1[1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U2 ( .A(MCInst_MC1_v3_3Inst_1_n3), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(MCInst_MC1_v3_3[1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .ZN(MCInst_MC1_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_0[2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_2_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_1[2]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_2[2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U2 ( .A(MCInst_MC1_v1_1Inst_2_n3), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_v1_1[2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U2 ( .A(MCInst_MC1_v1_2Inst_2_n3), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_v1_2[2]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U2 ( .A(MCInst_MC1_v2_1Inst_2_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_1[2]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U2 ( .A(MCInst_MC1_v2_2Inst_2_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_2[2]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC1_v2_3Inst_2_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(MCInst_MC1_v2_3[2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U2 ( .A(MCInst_MC1_v3_1Inst_2_n3), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(MCInst_MC1_v3_1[2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(MCInst_MC1_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC1_v3_3Inst_2_U1 ( .A(Red_MCInst_MC1_v3_3[2]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_v3_3[2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_3_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(MCInst_MC1_v0_1[3]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_3_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .Z(MCInst_MC1_v0_2[3]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_3_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        MCInst_MC1_v1_3[3]), .Z(MCInst_MC1_v1_1[3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U3 ( .A(MCInst_MC1_v1_2Inst_3_n6), .B(
        MCInst_MC1_v1_2Inst_3_n5), .ZN(MCInst_MC1_v1_2[3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U2 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC1_v1_2Inst_3_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .Z(MCInst_MC1_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC1_v2_1Inst_3_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(MCInst_MC1_v2_1[3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U2 ( .A(MCInst_MC1_v2_2Inst_3_n3), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(MCInst_MC1_v2_2[3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U2 ( .A(MCInst_MC1_v2_3Inst_3_n3), .B(
        MCInst_MC1_v2_0[3]), .ZN(MCInst_MC1_v2_3[3]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U1 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v2_0[2]), .ZN(MCInst_MC1_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC1_v3_1Inst_3_U1 ( .A(Red_MCInst_MC1_v3_3[2]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_v3_1[3]) );
  XOR2_X1 MCInst_MC1_v3_3Inst_3_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_v3_3[3]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_0_n8), .B(MCInst_MC1_r0Inst_XORInst_0_0_n7), .ZN(MC_output[56]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_2[1]), .B(
        MCInst_MC1_v1_0_0_), .ZN(MCInst_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_1_n8), .B(MCInst_MC1_r0Inst_XORInst_0_1_n7), .ZN(MC_output[57]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_0[1]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_0[1]), .B(
        MCInst_MC1_v3_0[1]), .Z(MCInst_MC1_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_2_n8), .B(MCInst_MC1_r0Inst_XORInst_0_2_n7), .ZN(MC_output[58]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_0[2]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r0Inst_XORInst_0_3_n8), .B(MCInst_MC1_r0Inst_XORInst_0_3_n7), .ZN(MC_output[59]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_0_n8), .B(MCInst_MC1_r1Inst_XORInst_0_0_n7), .ZN(MC_output[40]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_1[0]), .B(
        MCInst_MC1_v1_1[0]), .ZN(MCInst_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_1[0]), .Z(MCInst_MC1_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_1_n8), .B(MCInst_MC1_r1Inst_XORInst_0_1_n7), .ZN(MC_output[41]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v1_1[1]), .ZN(MCInst_MC1_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_1[1]), .B(
        MCInst_MC1_v3_1[1]), .Z(MCInst_MC1_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_2_n8), .B(MCInst_MC1_r1Inst_XORInst_0_2_n7), .ZN(MC_output[42]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_1[2]), .B(
        MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_1[2]), .B(
        MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r1Inst_XORInst_0_3_n8), .B(MCInst_MC1_r1Inst_XORInst_0_3_n7), .ZN(MC_output[43]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_1[3]), .B(
        MCInst_MC1_v1_1[3]), .ZN(MCInst_MC1_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_1[3]), .B(
        MCInst_MC1_v3_1[3]), .Z(MCInst_MC1_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_0_n8), .B(MCInst_MC1_r2Inst_XORInst_0_0_n7), .ZN(MC_output[24]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_2[0]), .B(
        MCInst_MC1_v1_2[0]), .ZN(MCInst_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC1_v0_2[0]), .B(
        MCInst_MC1_v3_2[0]), .Z(MCInst_MC1_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_1_n8), .B(MCInst_MC1_r2Inst_XORInst_0_1_n7), .ZN(MC_output[25]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_2[1]), .B(
        MCInst_MC1_v1_2[1]), .ZN(MCInst_MC1_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_2[1]), .B(
        MCInst_MC1_v3_0[3]), .Z(MCInst_MC1_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_2_n8), .B(MCInst_MC1_r2Inst_XORInst_0_2_n7), .ZN(MC_output[26]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_2[2]), .B(
        MCInst_MC1_v1_2[2]), .ZN(MCInst_MC1_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC1_v0_2[2]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(MCInst_MC1_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r2Inst_XORInst_0_3_n8), .B(MCInst_MC1_r2Inst_XORInst_0_3_n7), .ZN(MC_output[27]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_2[3]), .B(
        MCInst_MC1_v1_2[3]), .ZN(MCInst_MC1_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_2[3]), .B(
        MCInst_MC1_v3_2[3]), .Z(MCInst_MC1_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_0_n8), .B(MCInst_MC1_r3Inst_XORInst_0_0_n7), .ZN(MC_output[8]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC1_v2_3[0]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(MCInst_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_1[0]), .B(
        MCInst_MC1_v3_3[0]), .Z(MCInst_MC1_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_1_n8), .B(MCInst_MC1_r3Inst_XORInst_0_1_n7), .ZN(MC_output[9]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC1_v2_3[1]), .B(
        MCInst_MC1_v1_3[1]), .ZN(MCInst_MC1_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC1_v0_3[1]), .B(
        MCInst_MC1_v3_3[1]), .Z(MCInst_MC1_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_2_n8), .B(MCInst_MC1_r3Inst_XORInst_0_2_n7), .ZN(MC_output[10]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC1_v2_3[2]), .B(
        MCInst_MC1_v1_3[2]), .ZN(MCInst_MC1_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        MCInst_MC1_v3_3[2]), .Z(MCInst_MC1_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC1_r3Inst_XORInst_0_3_n8), .B(MCInst_MC1_r3Inst_XORInst_0_3_n7), .ZN(MC_output[11]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC1_v2_3[3]), .B(
        MCInst_MC1_v1_3[3]), .ZN(MCInst_MC1_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        MCInst_MC1_v3_3[3]), .Z(MCInst_MC1_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst_MC2_U2 ( .A(ShiftRowsOutput[20]), .Z(MCInst_MC2_v2_3[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U2 ( .A(MCInst_MC2_v0_2Inst_0_n3), .B(
        Red_MCInst_MC2_v0_1[0]), .ZN(MCInst_MC2_v0_2[0]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .ZN(MCInst_MC2_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v1_1Inst_0_U1 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .Z(MCInst_MC2_v1_1[0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U2 ( .A(MCInst_MC2_v1_2Inst_0_n3), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_v1_2[0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v2_1Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(MCInst_MC2_v2_1[0]) );
  XOR2_X1 MCInst_MC2_v2_2Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(MCInst_MC2_v2_2[0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U3 ( .A(MCInst_MC2_v2_3Inst_0_n6), .B(
        MCInst_MC2_v2_3Inst_0_n5), .ZN(MCInst_MC2_v2_3[0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC2_v2_3Inst_0_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC2_v3_1Inst_0_U1 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_v3_1[0]) );
  XOR2_X1 MCInst_MC2_v3_2Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_v3_2[0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U2 ( .A(MCInst_MC2_v3_3Inst_0_n3), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(MCInst_MC2_v3_3[0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(MCInst_MC2_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC2_v0_0Inst_1_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_0[1]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_1_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v0_3[3]), .Z(MCInst_MC2_v0_1[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U2 ( .A(MCInst_MC2_v0_2Inst_1_n3), .B(
        Red_MCInst_MC2_v0_1[0]), .ZN(MCInst_MC2_v0_2[1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .ZN(MCInst_MC2_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_3[1]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[3]), .Z(MCInst_MC2_v1_1[1]) );
  XOR2_X1 MCInst_MC2_v1_2Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .Z(MCInst_MC2_v1_2[1]) );
  XOR2_X1 MCInst_MC2_v1_3Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_1[2]), .Z(MCInst_MC2_v1_3[1]) );
  XOR2_X1 MCInst_MC2_v2_0Inst_1_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(MCInst_MC2_v2_0[1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U2 ( .A(MCInst_MC2_v2_1Inst_1_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_1[1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U3 ( .A(MCInst_MC2_v2_2Inst_1_n6), .B(
        MCInst_MC2_v2_2Inst_1_n5), .ZN(MCInst_MC2_v2_2[1]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC2_v2_2Inst_1_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC2_v3_0Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_v3_0[1]) );
  XOR2_X1 MCInst_MC2_v3_1Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_v3_1[1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U2 ( .A(MCInst_MC2_v3_3Inst_1_n3), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(MCInst_MC2_v3_3[1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .ZN(MCInst_MC2_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_0[2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_2_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_1[2]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_2[2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U2 ( .A(MCInst_MC2_v1_1Inst_2_n3), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_v1_1[2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U2 ( .A(MCInst_MC2_v1_2Inst_2_n3), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_v1_2[2]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U2 ( .A(MCInst_MC2_v2_1Inst_2_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_1[2]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U2 ( .A(MCInst_MC2_v2_2Inst_2_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_2[2]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC2_v2_3Inst_2_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(MCInst_MC2_v2_3[2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U2 ( .A(MCInst_MC2_v3_1Inst_2_n3), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(MCInst_MC2_v3_1[2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(MCInst_MC2_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC2_v3_3Inst_2_U1 ( .A(Red_MCInst_MC2_v3_3[2]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_v3_3[2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_3_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(MCInst_MC2_v0_1[3]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_3_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .Z(MCInst_MC2_v0_2[3]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_3_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        MCInst_MC2_v1_3[3]), .Z(MCInst_MC2_v1_1[3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U3 ( .A(MCInst_MC2_v1_2Inst_3_n6), .B(
        MCInst_MC2_v1_2Inst_3_n5), .ZN(MCInst_MC2_v1_2[3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U2 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC2_v1_2Inst_3_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .Z(MCInst_MC2_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC2_v2_1Inst_3_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(MCInst_MC2_v2_1[3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U2 ( .A(MCInst_MC2_v2_2Inst_3_n3), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(MCInst_MC2_v2_2[3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U2 ( .A(MCInst_MC2_v2_3Inst_3_n3), .B(
        MCInst_MC2_v2_0[3]), .ZN(MCInst_MC2_v2_3[3]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U1 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v2_0[2]), .ZN(MCInst_MC2_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC2_v3_1Inst_3_U1 ( .A(Red_MCInst_MC2_v3_3[2]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_v3_1[3]) );
  XOR2_X1 MCInst_MC2_v3_3Inst_3_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_v3_3[3]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_0_n8), .B(MCInst_MC2_r0Inst_XORInst_0_0_n7), .ZN(MC_output[52]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_2[1]), .B(
        MCInst_MC2_v1_0_0_), .ZN(MCInst_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_1_n8), .B(MCInst_MC2_r0Inst_XORInst_0_1_n7), .ZN(MC_output[53]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_0[1]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_0[1]), .B(
        MCInst_MC2_v3_0[1]), .Z(MCInst_MC2_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_2_n8), .B(MCInst_MC2_r0Inst_XORInst_0_2_n7), .ZN(MC_output[54]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_0[2]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r0Inst_XORInst_0_3_n8), .B(MCInst_MC2_r0Inst_XORInst_0_3_n7), .ZN(MC_output[55]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_0_n8), .B(MCInst_MC2_r1Inst_XORInst_0_0_n7), .ZN(MC_output[36]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_1[0]), .B(
        MCInst_MC2_v1_1[0]), .ZN(MCInst_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_1[0]), .Z(MCInst_MC2_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_1_n8), .B(MCInst_MC2_r1Inst_XORInst_0_1_n7), .ZN(MC_output[37]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v1_1[1]), .ZN(MCInst_MC2_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_1[1]), .B(
        MCInst_MC2_v3_1[1]), .Z(MCInst_MC2_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_2_n8), .B(MCInst_MC2_r1Inst_XORInst_0_2_n7), .ZN(MC_output[38]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_1[2]), .B(
        MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_1[2]), .B(
        MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r1Inst_XORInst_0_3_n8), .B(MCInst_MC2_r1Inst_XORInst_0_3_n7), .ZN(MC_output[39]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_1[3]), .B(
        MCInst_MC2_v1_1[3]), .ZN(MCInst_MC2_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_1[3]), .B(
        MCInst_MC2_v3_1[3]), .Z(MCInst_MC2_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_0_n8), .B(MCInst_MC2_r2Inst_XORInst_0_0_n7), .ZN(MC_output[20]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_2[0]), .B(
        MCInst_MC2_v1_2[0]), .ZN(MCInst_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC2_v0_2[0]), .B(
        MCInst_MC2_v3_2[0]), .Z(MCInst_MC2_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_1_n8), .B(MCInst_MC2_r2Inst_XORInst_0_1_n7), .ZN(MC_output[21]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_2[1]), .B(
        MCInst_MC2_v1_2[1]), .ZN(MCInst_MC2_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_2[1]), .B(
        MCInst_MC2_v3_0[3]), .Z(MCInst_MC2_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_2_n8), .B(MCInst_MC2_r2Inst_XORInst_0_2_n7), .ZN(MC_output[22]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_2[2]), .B(
        MCInst_MC2_v1_2[2]), .ZN(MCInst_MC2_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC2_v0_2[2]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(MCInst_MC2_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r2Inst_XORInst_0_3_n8), .B(MCInst_MC2_r2Inst_XORInst_0_3_n7), .ZN(MC_output[23]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_2[3]), .B(
        MCInst_MC2_v1_2[3]), .ZN(MCInst_MC2_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_2[3]), .B(
        MCInst_MC2_v3_2[3]), .Z(MCInst_MC2_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_0_n8), .B(MCInst_MC2_r3Inst_XORInst_0_0_n7), .ZN(MC_output[4]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC2_v2_3[0]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(MCInst_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_1[0]), .B(
        MCInst_MC2_v3_3[0]), .Z(MCInst_MC2_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_1_n8), .B(MCInst_MC2_r3Inst_XORInst_0_1_n7), .ZN(MC_output[5]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC2_v2_3[1]), .B(
        MCInst_MC2_v1_3[1]), .ZN(MCInst_MC2_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC2_v0_3[1]), .B(
        MCInst_MC2_v3_3[1]), .Z(MCInst_MC2_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_2_n8), .B(MCInst_MC2_r3Inst_XORInst_0_2_n7), .ZN(MC_output[6]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC2_v2_3[2]), .B(
        MCInst_MC2_v1_3[2]), .ZN(MCInst_MC2_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        MCInst_MC2_v3_3[2]), .Z(MCInst_MC2_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC2_r3Inst_XORInst_0_3_n8), .B(MCInst_MC2_r3Inst_XORInst_0_3_n7), .ZN(MC_output[7]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC2_v2_3[3]), .B(
        MCInst_MC2_v1_3[3]), .ZN(MCInst_MC2_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        MCInst_MC2_v3_3[3]), .Z(MCInst_MC2_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst_MC3_U2 ( .A(ShiftRowsOutput[16]), .Z(MCInst_MC3_v2_3[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U2 ( .A(MCInst_MC3_v0_2Inst_0_n3), .B(
        Red_MCInst_MC3_v0_1[0]), .ZN(MCInst_MC3_v0_2[0]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .ZN(MCInst_MC3_v0_2Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v1_1Inst_0_U1 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .Z(MCInst_MC3_v1_1[0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U2 ( .A(MCInst_MC3_v1_2Inst_0_n3), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_v1_2[0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_v1_2Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v2_1Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(MCInst_MC3_v2_1[0]) );
  XOR2_X1 MCInst_MC3_v2_2Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(MCInst_MC3_v2_2[0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U3 ( .A(MCInst_MC3_v2_3Inst_0_n6), .B(
        MCInst_MC3_v2_3Inst_0_n5), .ZN(MCInst_MC3_v2_3[0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_3Inst_0_n5) );
  XOR2_X1 MCInst_MC3_v2_3Inst_0_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_3Inst_0_n6) );
  XOR2_X1 MCInst_MC3_v3_1Inst_0_U1 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_v3_1[0]) );
  XOR2_X1 MCInst_MC3_v3_2Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_v3_2[0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U2 ( .A(MCInst_MC3_v3_3Inst_0_n3), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(MCInst_MC3_v3_3[0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(MCInst_MC3_v3_3Inst_0_n3) );
  XOR2_X1 MCInst_MC3_v0_0Inst_1_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_0[1]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_1_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v0_3[3]), .Z(MCInst_MC3_v0_1[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U2 ( .A(MCInst_MC3_v0_2Inst_1_n3), .B(
        Red_MCInst_MC3_v0_1[0]), .ZN(MCInst_MC3_v0_2[1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .ZN(MCInst_MC3_v0_2Inst_1_n3) );
  XOR2_X1 MCInst_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_3[1]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[3]), .Z(MCInst_MC3_v1_1[1]) );
  XOR2_X1 MCInst_MC3_v1_2Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .Z(MCInst_MC3_v1_2[1]) );
  XOR2_X1 MCInst_MC3_v1_3Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_1[2]), .Z(MCInst_MC3_v1_3[1]) );
  XOR2_X1 MCInst_MC3_v2_0Inst_1_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(MCInst_MC3_v2_0[1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U2 ( .A(MCInst_MC3_v2_1Inst_1_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_1[1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U3 ( .A(MCInst_MC3_v2_2Inst_1_n6), .B(
        MCInst_MC3_v2_2Inst_1_n5), .ZN(MCInst_MC3_v2_2[1]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_2Inst_1_n5) );
  XOR2_X1 MCInst_MC3_v2_2Inst_1_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_2Inst_1_n6) );
  XOR2_X1 MCInst_MC3_v3_0Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_v3_0[1]) );
  XOR2_X1 MCInst_MC3_v3_1Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_v3_1[1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U2 ( .A(MCInst_MC3_v3_3Inst_1_n3), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(MCInst_MC3_v3_3[1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .ZN(MCInst_MC3_v3_3Inst_1_n3) );
  XOR2_X1 MCInst_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_0[2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_2_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_1[2]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_2[2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U2 ( .A(MCInst_MC3_v1_1Inst_2_n3), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_v1_1[2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U2 ( .A(MCInst_MC3_v1_2Inst_2_n3), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_v1_2[2]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U2 ( .A(MCInst_MC3_v2_1Inst_2_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_1[2]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U2 ( .A(MCInst_MC3_v2_2Inst_2_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_2[2]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_2Inst_2_n3) );
  XOR2_X1 MCInst_MC3_v2_3Inst_2_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(MCInst_MC3_v2_3[2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U2 ( .A(MCInst_MC3_v3_1Inst_2_n3), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(MCInst_MC3_v3_1[2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(MCInst_MC3_v3_1Inst_2_n3) );
  XOR2_X1 MCInst_MC3_v3_3Inst_2_U1 ( .A(Red_MCInst_MC3_v3_3[2]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_v3_3[2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_3_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(MCInst_MC3_v0_1[3]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_3_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .Z(MCInst_MC3_v0_2[3]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_3_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        MCInst_MC3_v1_3[3]), .Z(MCInst_MC3_v1_1[3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U3 ( .A(MCInst_MC3_v1_2Inst_3_n6), .B(
        MCInst_MC3_v1_2Inst_3_n5), .ZN(MCInst_MC3_v1_2[3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U2 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_v1_2Inst_3_n5) );
  XOR2_X1 MCInst_MC3_v1_2Inst_3_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .Z(MCInst_MC3_v1_2Inst_3_n6) );
  XOR2_X1 MCInst_MC3_v2_1Inst_3_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(MCInst_MC3_v2_1[3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U2 ( .A(MCInst_MC3_v2_2Inst_3_n3), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(MCInst_MC3_v2_2[3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U2 ( .A(MCInst_MC3_v2_3Inst_3_n3), .B(
        MCInst_MC3_v2_0[3]), .ZN(MCInst_MC3_v2_3[3]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U1 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v2_0[2]), .ZN(MCInst_MC3_v2_3Inst_3_n3) );
  XOR2_X1 MCInst_MC3_v3_1Inst_3_U1 ( .A(Red_MCInst_MC3_v3_3[2]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_v3_1[3]) );
  XOR2_X1 MCInst_MC3_v3_3Inst_3_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_v3_3[3]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_0_n8), .B(MCInst_MC3_r0Inst_XORInst_0_0_n7), .ZN(MC_output[48]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_2[1]), .B(
        MCInst_MC3_v1_0_0_), .ZN(MCInst_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_1_n8), .B(MCInst_MC3_r0Inst_XORInst_0_1_n7), .ZN(MC_output[49]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_0[1]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_0[1]), .B(
        MCInst_MC3_v3_0[1]), .Z(MCInst_MC3_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_2_n8), .B(MCInst_MC3_r0Inst_XORInst_0_2_n7), .ZN(MC_output[50]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_0[2]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r0Inst_XORInst_0_3_n8), .B(MCInst_MC3_r0Inst_XORInst_0_3_n7), .ZN(MC_output[51]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_0_n8), .B(MCInst_MC3_r1Inst_XORInst_0_0_n7), .ZN(MC_output[32]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_1[0]), .B(
        MCInst_MC3_v1_1[0]), .ZN(MCInst_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_1[0]), .Z(MCInst_MC3_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_1_n8), .B(MCInst_MC3_r1Inst_XORInst_0_1_n7), .ZN(MC_output[33]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v1_1[1]), .ZN(MCInst_MC3_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_1[1]), .B(
        MCInst_MC3_v3_1[1]), .Z(MCInst_MC3_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_2_n8), .B(MCInst_MC3_r1Inst_XORInst_0_2_n7), .ZN(MC_output[34]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_1[2]), .B(
        MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_1[2]), .B(
        MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r1Inst_XORInst_0_3_n8), .B(MCInst_MC3_r1Inst_XORInst_0_3_n7), .ZN(MC_output[35]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_1[3]), .B(
        MCInst_MC3_v1_1[3]), .ZN(MCInst_MC3_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_1[3]), .B(
        MCInst_MC3_v3_1[3]), .Z(MCInst_MC3_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_0_n8), .B(MCInst_MC3_r2Inst_XORInst_0_0_n7), .ZN(MC_output[16]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_2[0]), .B(
        MCInst_MC3_v1_2[0]), .ZN(MCInst_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U1 ( .A(MCInst_MC3_v0_2[0]), .B(
        MCInst_MC3_v3_2[0]), .Z(MCInst_MC3_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_1_n8), .B(MCInst_MC3_r2Inst_XORInst_0_1_n7), .ZN(MC_output[17]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_2[1]), .B(
        MCInst_MC3_v1_2[1]), .ZN(MCInst_MC3_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_2[1]), .B(
        MCInst_MC3_v3_0[3]), .Z(MCInst_MC3_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_2_n8), .B(MCInst_MC3_r2Inst_XORInst_0_2_n7), .ZN(MC_output[18]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_2[2]), .B(
        MCInst_MC3_v1_2[2]), .ZN(MCInst_MC3_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U1 ( .A(MCInst_MC3_v0_2[2]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(MCInst_MC3_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r2Inst_XORInst_0_3_n8), .B(MCInst_MC3_r2Inst_XORInst_0_3_n7), .ZN(MC_output[19]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_2[3]), .B(
        MCInst_MC3_v1_2[3]), .ZN(MCInst_MC3_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_2[3]), .B(
        MCInst_MC3_v3_2[3]), .Z(MCInst_MC3_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_0_n8), .B(MCInst_MC3_r3Inst_XORInst_0_0_n7), .ZN(MC_output[0]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U2 ( .A(MCInst_MC3_v2_3[0]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(MCInst_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_1[0]), .B(
        MCInst_MC3_v3_3[0]), .Z(MCInst_MC3_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_1_n8), .B(MCInst_MC3_r3Inst_XORInst_0_1_n7), .ZN(MC_output[1]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U2 ( .A(MCInst_MC3_v2_3[1]), .B(
        MCInst_MC3_v1_3[1]), .ZN(MCInst_MC3_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U1 ( .A(MCInst_MC3_v0_3[1]), .B(
        MCInst_MC3_v3_3[1]), .Z(MCInst_MC3_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_2_n8), .B(MCInst_MC3_r3Inst_XORInst_0_2_n7), .ZN(MC_output[2]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U2 ( .A(MCInst_MC3_v2_3[2]), .B(
        MCInst_MC3_v1_3[2]), .ZN(MCInst_MC3_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        MCInst_MC3_v3_3[2]), .Z(MCInst_MC3_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst_MC3_r3Inst_XORInst_0_3_n8), .B(MCInst_MC3_r3Inst_XORInst_0_3_n7), .ZN(MC_output[3]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U2 ( .A(MCInst_MC3_v2_3[3]), .B(
        MCInst_MC3_v1_3[3]), .ZN(MCInst_MC3_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        MCInst_MC3_v3_3[3]), .Z(MCInst_MC3_r3Inst_XORInst_0_3_n8) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(MC_output[0]), .CK(clk), .Q(
        SubCellInput2[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(MC_output[1]), .CK(clk), .Q(
        SubCellInput2[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(MC_output[2]), .CK(clk), .Q(
        SubCellInput2[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(MC_output[3]), .CK(clk), .Q(
        SubCellInput2[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(MC_output[4]), .CK(clk), .Q(
        SubCellInput2[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(MC_output[5]), .CK(clk), .Q(
        SubCellInput2[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(MC_output[6]), .CK(clk), .Q(
        SubCellInput2[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(MC_output[7]), .CK(clk), .Q(
        SubCellInput2[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(MC_output[8]), .CK(clk), .Q(
        SubCellInput2[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(MC_output[9]), .CK(clk), .Q(
        SubCellInput2[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(MC_output[10]), .CK(clk), .Q(
        SubCellInput2[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(MC_output[11]), .CK(clk), .Q(
        SubCellInput2[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(MC_output[12]), .CK(clk), .Q(
        SubCellInput2[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(MC_output[13]), .CK(clk), .Q(
        SubCellInput2[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(MC_output[14]), .CK(clk), .Q(
        SubCellInput2[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(MC_output[15]), .CK(clk), .Q(
        SubCellInput2[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(MC_output[16]), .CK(clk), .Q(
        SubCellInput2[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(MC_output[17]), .CK(clk), .Q(
        SubCellInput2[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(MC_output[18]), .CK(clk), .Q(
        SubCellInput2[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(MC_output[19]), .CK(clk), .Q(
        SubCellInput2[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(MC_output[20]), .CK(clk), .Q(
        SubCellInput2[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(MC_output[21]), .CK(clk), .Q(
        SubCellInput2[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(MC_output[22]), .CK(clk), .Q(
        SubCellInput2[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(MC_output[23]), .CK(clk), .Q(
        SubCellInput2[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(MC_output[24]), .CK(clk), .Q(
        SubCellInput2[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(MC_output[25]), .CK(clk), .Q(
        SubCellInput2[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(MC_output[26]), .CK(clk), .Q(
        SubCellInput2[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(MC_output[27]), .CK(clk), .Q(
        SubCellInput2[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(MC_output[28]), .CK(clk), .Q(
        SubCellInput2[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(MC_output[29]), .CK(clk), .Q(
        SubCellInput2[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(MC_output[30]), .CK(clk), .Q(
        SubCellInput2[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(MC_output[31]), .CK(clk), .Q(
        SubCellInput2[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(MC_output[32]), .CK(clk), .Q(
        SubCellInput2[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(MC_output[33]), .CK(clk), .Q(
        SubCellInput2[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(MC_output[34]), .CK(clk), .Q(
        SubCellInput2[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(MC_output[35]), .CK(clk), .Q(
        SubCellInput2[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(MC_output[36]), .CK(clk), .Q(
        SubCellInput2[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(MC_output[37]), .CK(clk), .Q(
        SubCellInput2[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(MC_output[38]), .CK(clk), .Q(
        SubCellInput2[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(MC_output[39]), .CK(clk), .Q(
        SubCellInput2[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(MC_output[40]), .CK(clk), .Q(
        SubCellInput2[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(MC_output[41]), .CK(clk), .Q(
        SubCellInput2[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(MC_output[42]), .CK(clk), .Q(
        SubCellInput2[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(MC_output[43]), .CK(clk), .Q(
        SubCellInput2[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(MC_output[44]), .CK(clk), .Q(
        SubCellInput2[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(MC_output[45]), .CK(clk), .Q(
        SubCellInput2[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(MC_output[46]), .CK(clk), .Q(
        SubCellInput2[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(MC_output[47]), .CK(clk), .Q(
        SubCellInput2[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(MC_output[48]), .CK(clk), .Q(
        SubCellInput2[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(MC_output[49]), .CK(clk), .Q(
        SubCellInput2[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(MC_output[50]), .CK(clk), .Q(
        SubCellInput2[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(MC_output[51]), .CK(clk), .Q(
        SubCellInput2[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(MC_output[52]), .CK(clk), .Q(
        SubCellInput2[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(MC_output[53]), .CK(clk), .Q(
        SubCellInput2[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(MC_output[54]), .CK(clk), .Q(
        SubCellInput2[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(MC_output[55]), .CK(clk), .Q(
        SubCellInput2[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(MC_output[56]), .CK(clk), .Q(
        SubCellInput2[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(MC_output[57]), .CK(clk), .Q(
        SubCellInput2[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(MC_output[58]), .CK(clk), .Q(
        SubCellInput2[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(MC_output[59]), .CK(clk), .Q(
        SubCellInput2[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(MC_output[60]), .CK(clk), .Q(
        SubCellInput2[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(MC_output[61]), .CK(clk), .Q(
        SubCellInput2[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(MC_output[62]), .CK(clk), .Q(
        SubCellInput2[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(MC_output[63]), .CK(clk), .Q(
        SubCellInput2[63]), .QN() );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_0_U5 ( .A1(SubCellInput2[2]), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_0_U4 ( .A(SubCellInput2[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U3 ( .A(SubCellInput2[0]), .B(
        SubCellInput2[3]), .Z(SubCellInst2_LFInst_0_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_0_LFInst_0_n8), .ZN(MCInst2_MC0_v3_2[3]) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_0_LFInst_0_n7), .B(
        SubCellInst2_LFInst_0_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_0_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_1_U9 ( .A1(SubCellInput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_1_U8 ( .A(SubCellInput2[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n21), .A2(SubCellInput2[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U5 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U3 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_1_U2 ( .A(SubCellInput2[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n19) );
  NAND2_X2 SubCellInst2_LFInst_0_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n25), .ZN(Red_MCInst2_MC0_v3_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n28), .ZN(MCInst2_MC0_v3_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_2_U6 ( .A(SubCellInput2[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_0_LFInst_2_n25), .B(SubCellInput2[2]), .Z(
        SubCellInst2_LFInst_0_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U4 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n23), .A2(SubCellInput2[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_0_LFInst_2_n22), .B(SubCellInput2[1]), .Z(
        SubCellInst2_LFInst_0_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_2_U1 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U9 ( .A1(SubCellInput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n23), .A2(SubCellInput2[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_3_U7 ( .A1(SubCellInput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U4 ( .A1(SubCellInput2[2]), .A2(
        SubCellInput2[0]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_3_U3 ( .A(SubCellInput2[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U2 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n25), .ZN(Red_MCInst2_MC0_v3_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_0_U5 ( .A1(SubCellInput2[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_0_U4 ( .A(SubCellInput2[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U3 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[7]), .Z(SubCellInst2_LFInst_1_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_1_LFInst_0_n8), .ZN(MCInst2_MC3_v3_2[3]) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_1_LFInst_0_n7), .B(
        SubCellInst2_LFInst_1_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_1_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_1_U9 ( .A1(SubCellInput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_1_U8 ( .A(SubCellInput2[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n21), .A2(SubCellInput2[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U5 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U3 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_1_U2 ( .A(SubCellInput2[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n19) );
  NAND2_X2 SubCellInst2_LFInst_1_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n25), .ZN(Red_MCInst2_MC3_v3_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U9 ( .A1(SubCellInput2[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U8 ( .A1(SubCellInput2[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_2_U7 ( .A(SubCellInput2[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_1_LFInst_2_n23), .B(SubCellInput2[6]), .Z(
        SubCellInst2_LFInst_1_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U4 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n22), .A2(SubCellInput2[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U2 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n28), .ZN(MCInst2_MC3_v3_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U9 ( .A1(SubCellInput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n23), .A2(SubCellInput2[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_3_U7 ( .A1(SubCellInput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U4 ( .A1(SubCellInput2[6]), .A2(
        SubCellInput2[4]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_3_U3 ( .A(SubCellInput2[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U2 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n25), .ZN(Red_MCInst2_MC3_v3_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_0_U5 ( .A1(SubCellInput2[10]), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_0_U4 ( .A(SubCellInput2[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U3 ( .A(SubCellInput2[8]), .B(
        SubCellInput2[11]), .Z(SubCellInst2_LFInst_2_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_2_LFInst_0_n8), .ZN(MCInst2_MC2_v3_2[3]) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_2_LFInst_0_n7), .B(
        SubCellInst2_LFInst_2_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_2_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_1_U9 ( .A1(SubCellInput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_1_U8 ( .A(SubCellInput2[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n21), .A2(SubCellInput2[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U5 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U3 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_1_U2 ( .A(SubCellInput2[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n19) );
  NAND2_X2 SubCellInst2_LFInst_2_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n25), .ZN(Red_MCInst2_MC2_v3_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n28), .ZN(MCInst2_MC2_v3_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_2_U6 ( .A(SubCellInput2[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_2_LFInst_2_n25), .B(SubCellInput2[10]), .Z(
        SubCellInst2_LFInst_2_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U4 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n23), .A2(SubCellInput2[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_2_LFInst_2_n22), .B(SubCellInput2[9]), .Z(
        SubCellInst2_LFInst_2_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_2_U1 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U9 ( .A1(SubCellInput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n23), .A2(SubCellInput2[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_3_U7 ( .A1(SubCellInput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U4 ( .A1(SubCellInput2[10]), .A2(
        SubCellInput2[8]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_3_U3 ( .A(SubCellInput2[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U2 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n25), .ZN(Red_MCInst2_MC2_v3_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_0_U5 ( .A1(SubCellInput2[14]), .A2(
        SubCellInst2_LFInst_3_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_0_U4 ( .A(SubCellInput2[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U3 ( .A(SubCellInput2[12]), .B(
        SubCellInput2[15]), .Z(SubCellInst2_LFInst_3_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_3_LFInst_0_n8), .ZN(MCInst2_MC1_v3_2[3]) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_3_LFInst_0_n7), .B(
        SubCellInst2_LFInst_3_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_3_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_1_U9 ( .A1(SubCellInput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_1_U8 ( .A(SubCellInput2[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n21), .A2(SubCellInput2[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U5 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U3 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_1_U2 ( .A(SubCellInput2[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n19) );
  NAND2_X2 SubCellInst2_LFInst_3_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n25), .ZN(Red_MCInst2_MC1_v3_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n28), .ZN(MCInst2_MC1_v3_0[3]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_2_U6 ( .A(SubCellInput2[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_3_LFInst_2_n25), .B(SubCellInput2[14]), .Z(
        SubCellInst2_LFInst_3_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U4 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n23), .A2(SubCellInput2[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_3_LFInst_2_n22), .B(SubCellInput2[13]), .Z(
        SubCellInst2_LFInst_3_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_2_U1 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U9 ( .A1(SubCellInput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n23), .A2(SubCellInput2[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_3_U7 ( .A1(SubCellInput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U4 ( .A1(SubCellInput2[14]), .A2(
        SubCellInput2[12]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_3_U3 ( .A(SubCellInput2[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U2 ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n25), .ZN(Red_MCInst2_MC1_v3_1[2]) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U4 ( .A(
        SubCellInst2_LFInst_4_LFInst_0_n6), .B(
        SubCellInst2_LFInst_4_LFInst_0_n5), .ZN(ShiftRowsOutput2[24]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_0_U3 ( .A1(SubCellInput2[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_0_n4), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n5) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_0_U2 ( .A(SubCellInput2[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n4) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U1 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[19]), .Z(SubCellInst2_LFInst_4_LFInst_0_n6) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_1_U9 ( .A1(SubCellInput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_1_U8 ( .A(SubCellInput2[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n21), .A2(SubCellInput2[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U5 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U3 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_1_U2 ( .A(SubCellInput2[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n25), .ZN(MCInst2_MC1_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U9 ( .A1(SubCellInput2[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U8 ( .A1(SubCellInput2[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_2_U7 ( .A(SubCellInput2[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_4_LFInst_2_n23), .B(SubCellInput2[18]), .Z(
        SubCellInst2_LFInst_4_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U4 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n22), .A2(SubCellInput2[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U2 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n22) );
  NAND2_X2 SubCellInst2_LFInst_4_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n28), .ZN(MCInst2_MC1_v2_0[3]) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n25), .A2(SubCellInput2[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n25), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n23), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n24) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n22), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n23) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U6 ( .A1(SubCellInput2[18]), .A2(
        SubCellInput2[16]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n21) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_3_U5 ( .A(SubCellInput2[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U4 ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n25) );
  AND2_X1 SubCellInst2_LFInst_4_LFInst_3_U3 ( .A1(SubCellInput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n26), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U2 ( .A1(SubCellInput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n19) );
  OR2_X2 SubCellInst2_LFInst_4_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n19), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n20), .ZN(Red_MCInst2_MC1_v2_2[1]) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U4 ( .A(
        SubCellInst2_LFInst_5_LFInst_0_n6), .B(
        SubCellInst2_LFInst_5_LFInst_0_n5), .ZN(ShiftRowsOutput2[28]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_0_U3 ( .A1(SubCellInput2[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_0_n4), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n5) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_0_U2 ( .A(SubCellInput2[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n4) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U1 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[23]), .Z(SubCellInst2_LFInst_5_LFInst_0_n6) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_1_U9 ( .A1(SubCellInput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_1_U8 ( .A(SubCellInput2[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n21), .A2(SubCellInput2[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U5 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U3 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_1_U2 ( .A(SubCellInput2[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n25), .ZN(MCInst2_MC0_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U9 ( .A1(SubCellInput2[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U8 ( .A1(SubCellInput2[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_2_U7 ( .A(SubCellInput2[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_5_LFInst_2_n23), .B(SubCellInput2[22]), .Z(
        SubCellInst2_LFInst_5_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U4 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n22), .A2(SubCellInput2[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U2 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n22) );
  NAND2_X2 SubCellInst2_LFInst_5_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n28), .ZN(MCInst2_MC0_v2_0[3]) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n25), .A2(SubCellInput2[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n25), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n23), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n24) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n22), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n23) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U6 ( .A1(SubCellInput2[22]), .A2(
        SubCellInput2[20]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n21) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_3_U5 ( .A(SubCellInput2[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U4 ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n25) );
  AND2_X1 SubCellInst2_LFInst_5_LFInst_3_U3 ( .A1(SubCellInput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n26), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U2 ( .A1(SubCellInput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n19) );
  OR2_X2 SubCellInst2_LFInst_5_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n19), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n20), .ZN(Red_MCInst2_MC0_v2_2[1]) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U4 ( .A(
        SubCellInst2_LFInst_6_LFInst_0_n6), .B(
        SubCellInst2_LFInst_6_LFInst_0_n5), .ZN(ShiftRowsOutput2[16]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_0_U3 ( .A1(SubCellInput2[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_0_n4), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n5) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_0_U2 ( .A(SubCellInput2[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n4) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U1 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[27]), .Z(SubCellInst2_LFInst_6_LFInst_0_n6) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_1_U9 ( .A1(SubCellInput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_1_U8 ( .A(SubCellInput2[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n21), .A2(SubCellInput2[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U5 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U3 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_1_U2 ( .A(SubCellInput2[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n25), .ZN(MCInst2_MC3_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U9 ( .A1(SubCellInput2[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U8 ( .A1(SubCellInput2[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_2_U7 ( .A(SubCellInput2[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_6_LFInst_2_n23), .B(SubCellInput2[26]), .Z(
        SubCellInst2_LFInst_6_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U4 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n22), .A2(SubCellInput2[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U2 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n22) );
  NAND2_X2 SubCellInst2_LFInst_6_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n28), .ZN(MCInst2_MC3_v2_0[3]) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n25), .A2(SubCellInput2[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n25), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n23), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n24) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n22), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n23) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U6 ( .A1(SubCellInput2[26]), .A2(
        SubCellInput2[24]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n21) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_3_U5 ( .A(SubCellInput2[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U4 ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n25) );
  AND2_X1 SubCellInst2_LFInst_6_LFInst_3_U3 ( .A1(SubCellInput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n26), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U2 ( .A1(SubCellInput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n19) );
  OR2_X2 SubCellInst2_LFInst_6_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n19), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n20), .ZN(Red_MCInst2_MC3_v2_2[1]) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U4 ( .A(
        SubCellInst2_LFInst_7_LFInst_0_n6), .B(
        SubCellInst2_LFInst_7_LFInst_0_n5), .ZN(ShiftRowsOutput2[20]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_0_U3 ( .A1(SubCellInput2[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_0_n4), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n5) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_0_U2 ( .A(SubCellInput2[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n4) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U1 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[31]), .Z(SubCellInst2_LFInst_7_LFInst_0_n6) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_1_U9 ( .A1(SubCellInput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_1_U8 ( .A(SubCellInput2[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n21), .A2(SubCellInput2[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U5 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U3 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_1_U2 ( .A(SubCellInput2[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n25), .ZN(MCInst2_MC2_v2_0[2]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U9 ( .A1(SubCellInput2[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U8 ( .A1(SubCellInput2[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_2_U7 ( .A(SubCellInput2[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_7_LFInst_2_n23), .B(SubCellInput2[30]), .Z(
        SubCellInst2_LFInst_7_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U4 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n22), .A2(SubCellInput2[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U2 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n22) );
  NAND2_X2 SubCellInst2_LFInst_7_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n28), .ZN(MCInst2_MC2_v2_0[3]) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U9 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n25), .A2(SubCellInput2[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n25), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n23), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n24) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U7 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n22), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n23) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U6 ( .A1(SubCellInput2[30]), .A2(
        SubCellInput2[28]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n21) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_3_U5 ( .A(SubCellInput2[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U4 ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n25) );
  AND2_X1 SubCellInst2_LFInst_7_LFInst_3_U3 ( .A1(SubCellInput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n26), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U2 ( .A1(SubCellInput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n19) );
  OR2_X2 SubCellInst2_LFInst_7_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n19), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n20), .ZN(Red_MCInst2_MC2_v2_2[1]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_0_U5 ( .A1(SubCellInput2[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_0_n7), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n8) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_0_U4 ( .A(SubCellInput2[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n7) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U3 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[35]), .Z(SubCellInst2_LFInst_8_LFInst_0_n9) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_8_LFInst_0_n10), .ZN(MCInst2_MC2_v1_0_0_) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_8_LFInst_0_n9), .B(
        SubCellInst2_LFInst_8_LFInst_0_n8), .Z(
        SubCellInst2_LFInst_8_LFInst_0_n10) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n25), .ZN(MCInst2_MC2_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_1_U8 ( .A1(SubCellInput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_1_U7 ( .A(SubCellInput2[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n21), .A2(SubCellInput2[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U4 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U2 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_1_U1 ( .A(SubCellInput2[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U9 ( .A1(SubCellInput2[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U8 ( .A1(SubCellInput2[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_2_U7 ( .A(SubCellInput2[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_8_LFInst_2_n23), .B(SubCellInput2[34]), .Z(
        SubCellInst2_LFInst_8_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U4 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n22), .A2(SubCellInput2[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U2 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n28), .ZN(MCInst2_MC2_v1_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U9 ( .A1(SubCellInput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n23), .A2(SubCellInput2[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_3_U7 ( .A1(SubCellInput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U4 ( .A1(SubCellInput2[34]), .A2(
        SubCellInput2[32]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_3_U3 ( .A(SubCellInput2[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U2 ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n25), .ZN(Red_MCInst2_MC2_v1_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_0_U5 ( .A1(SubCellInput2[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_0_n7), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n8) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_0_U4 ( .A(SubCellInput2[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n7) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U3 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[39]), .Z(SubCellInst2_LFInst_9_LFInst_0_n9) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_9_LFInst_0_n10), .ZN(MCInst2_MC1_v1_0_0_) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_9_LFInst_0_n9), .B(
        SubCellInst2_LFInst_9_LFInst_0_n8), .Z(
        SubCellInst2_LFInst_9_LFInst_0_n10) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n25), .ZN(MCInst2_MC1_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_1_U8 ( .A1(SubCellInput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_1_U7 ( .A(SubCellInput2[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n21), .A2(SubCellInput2[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U4 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U2 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_1_U1 ( .A(SubCellInput2[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U9 ( .A1(SubCellInput2[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U8 ( .A1(SubCellInput2[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_2_U7 ( .A(SubCellInput2[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_9_LFInst_2_n23), .B(SubCellInput2[38]), .Z(
        SubCellInst2_LFInst_9_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U4 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n22), .A2(SubCellInput2[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U2 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n28), .ZN(MCInst2_MC1_v1_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U9 ( .A1(SubCellInput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n23), .A2(SubCellInput2[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_3_U7 ( .A1(SubCellInput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U4 ( .A1(SubCellInput2[38]), .A2(
        SubCellInput2[36]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_3_U3 ( .A(SubCellInput2[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U2 ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n25), .ZN(Red_MCInst2_MC1_v1_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_0_U5 ( .A1(SubCellInput2[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_0_n7), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n8) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_0_U4 ( .A(SubCellInput2[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n7) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U3 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[43]), .Z(SubCellInst2_LFInst_10_LFInst_0_n9) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_10_LFInst_0_n10), .ZN(MCInst2_MC0_v1_0_0_) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_10_LFInst_0_n9), .B(
        SubCellInst2_LFInst_10_LFInst_0_n8), .Z(
        SubCellInst2_LFInst_10_LFInst_0_n10) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n25), .ZN(MCInst2_MC0_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_1_U8 ( .A1(SubCellInput2[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_1_U7 ( .A(SubCellInput2[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n21), .A2(SubCellInput2[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U4 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U2 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_1_U1 ( .A(SubCellInput2[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U9 ( .A1(SubCellInput2[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U8 ( .A1(SubCellInput2[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_2_U7 ( .A(SubCellInput2[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_10_LFInst_2_n23), .B(SubCellInput2[42]), .Z(
        SubCellInst2_LFInst_10_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U4 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n22), .A2(SubCellInput2[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U2 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n28), .ZN(MCInst2_MC0_v1_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U9 ( .A1(SubCellInput2[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n23), .A2(SubCellInput2[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_3_U7 ( .A1(SubCellInput2[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U4 ( .A1(SubCellInput2[42]), .A2(
        SubCellInput2[40]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_3_U3 ( .A(SubCellInput2[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U2 ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n25), .ZN(Red_MCInst2_MC0_v1_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_0_U5 ( .A1(SubCellInput2[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_0_n7), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n8) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_0_U4 ( .A(SubCellInput2[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n7) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U3 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[47]), .Z(SubCellInst2_LFInst_11_LFInst_0_n9) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_11_LFInst_0_n10), .ZN(MCInst2_MC3_v1_0_0_) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_11_LFInst_0_n9), .B(
        SubCellInst2_LFInst_11_LFInst_0_n8), .Z(
        SubCellInst2_LFInst_11_LFInst_0_n10) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n25), .ZN(MCInst2_MC3_v1_3[2]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U9 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_1_U8 ( .A1(SubCellInput2[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_1_U7 ( .A(SubCellInput2[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n21), .A2(SubCellInput2[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U5 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U4 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U3 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U2 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_1_U1 ( .A(SubCellInput2[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U8 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n24), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n28), .ZN(MCInst2_MC3_v1_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U7 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n26), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n28) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_2_U6 ( .A(SubCellInput2[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n27) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_11_LFInst_2_n25), .B(SubCellInput2[46]), .Z(
        SubCellInst2_LFInst_11_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U4 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n25) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n23), .A2(SubCellInput2[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n24) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U2 ( .A(
        SubCellInst2_LFInst_11_LFInst_2_n22), .B(SubCellInput2[45]), .Z(
        SubCellInst2_LFInst_11_LFInst_2_n23) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_2_U1 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U9 ( .A1(SubCellInput2[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n23), .A2(SubCellInput2[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_3_U7 ( .A1(SubCellInput2[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U4 ( .A1(SubCellInput2[46]), .A2(
        SubCellInput2[44]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_3_U3 ( .A(SubCellInput2[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U2 ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n25), .ZN(Red_MCInst2_MC3_v1_1[2]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_0_U5 ( .A1(SubCellInput2[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_0_U4 ( .A(SubCellInput2[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U3 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[51]), .Z(SubCellInst2_LFInst_12_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_12_LFInst_0_n8), .ZN(Red_MCInst2_MC3_v0_0[0]) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_12_LFInst_0_n7), .B(
        SubCellInst2_LFInst_12_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_12_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_1_U9 ( .A1(SubCellInput2[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_1_U8 ( .A(SubCellInput2[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n21), .A2(SubCellInput2[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U5 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U3 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_1_U2 ( .A(SubCellInput2[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n25), .ZN(Red_MCInst2_MC3_v0_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U9 ( .A1(SubCellInput2[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U8 ( .A1(SubCellInput2[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_2_U7 ( .A(SubCellInput2[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_12_LFInst_2_n23), .B(SubCellInput2[50]), .Z(
        SubCellInst2_LFInst_12_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U4 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n22), .A2(SubCellInput2[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U2 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n28), .ZN(MCInst2_MC3_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U9 ( .A1(SubCellInput2[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n23), .A2(SubCellInput2[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_3_U7 ( .A1(SubCellInput2[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U4 ( .A1(SubCellInput2[50]), .A2(
        SubCellInput2[48]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_3_U3 ( .A(SubCellInput2[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U2 ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n25), .ZN(Red_MCInst2_MC3_v0_1[0]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_0_U5 ( .A1(SubCellInput2[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_0_U4 ( .A(SubCellInput2[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U3 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[55]), .Z(SubCellInst2_LFInst_13_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_13_LFInst_0_n8), .ZN(Red_MCInst2_MC2_v0_0[0]) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_13_LFInst_0_n7), .B(
        SubCellInst2_LFInst_13_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_13_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_1_U9 ( .A1(SubCellInput2[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_1_U8 ( .A(SubCellInput2[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n21), .A2(SubCellInput2[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U5 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U3 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_1_U2 ( .A(SubCellInput2[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n25), .ZN(Red_MCInst2_MC2_v0_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U9 ( .A1(SubCellInput2[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U8 ( .A1(SubCellInput2[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_2_U7 ( .A(SubCellInput2[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_13_LFInst_2_n23), .B(SubCellInput2[54]), .Z(
        SubCellInst2_LFInst_13_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U4 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n22), .A2(SubCellInput2[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U2 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n28), .ZN(MCInst2_MC2_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U9 ( .A1(SubCellInput2[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n23), .A2(SubCellInput2[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_3_U7 ( .A1(SubCellInput2[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U4 ( .A1(SubCellInput2[54]), .A2(
        SubCellInput2[52]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_3_U3 ( .A(SubCellInput2[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U2 ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n25), .ZN(Red_MCInst2_MC2_v0_1[0]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_0_U5 ( .A1(SubCellInput2[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_0_U4 ( .A(SubCellInput2[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U3 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[59]), .Z(SubCellInst2_LFInst_14_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_14_LFInst_0_n8), .ZN(Red_MCInst2_MC1_v0_0[0]) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_14_LFInst_0_n7), .B(
        SubCellInst2_LFInst_14_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_14_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_1_U9 ( .A1(SubCellInput2[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_1_U8 ( .A(SubCellInput2[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n21), .A2(SubCellInput2[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U5 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U3 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_1_U2 ( .A(SubCellInput2[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n25), .ZN(Red_MCInst2_MC1_v0_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U9 ( .A1(SubCellInput2[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U8 ( .A1(SubCellInput2[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_2_U7 ( .A(SubCellInput2[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_14_LFInst_2_n23), .B(SubCellInput2[58]), .Z(
        SubCellInst2_LFInst_14_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U4 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n22), .A2(SubCellInput2[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U2 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n28), .ZN(MCInst2_MC1_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U9 ( .A1(SubCellInput2[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n23), .A2(SubCellInput2[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_3_U7 ( .A1(SubCellInput2[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U4 ( .A1(SubCellInput2[58]), .A2(
        SubCellInput2[56]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_3_U3 ( .A(SubCellInput2[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U2 ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n25), .ZN(Red_MCInst2_MC1_v0_1[0]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_0_U5 ( .A1(SubCellInput2[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_0_n5), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n6) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_0_U4 ( .A(SubCellInput2[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n5) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U3 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[63]), .Z(SubCellInst2_LFInst_15_LFInst_0_n7) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_0_U2 ( .A(
        SubCellInst2_LFInst_15_LFInst_0_n8), .ZN(Red_MCInst2_MC0_v0_0[0]) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U1 ( .A(
        SubCellInst2_LFInst_15_LFInst_0_n7), .B(
        SubCellInst2_LFInst_15_LFInst_0_n6), .Z(
        SubCellInst2_LFInst_15_LFInst_0_n8) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U10 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n24), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n25) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_1_U9 ( .A1(SubCellInput2[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n22), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n24) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_1_U8 ( .A(SubCellInput2[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n22) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U7 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n21), .A2(SubCellInput2[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n26) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n20), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n23), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n21) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U5 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n23) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n19), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n18), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n20) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U3 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n18) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_1_U2 ( .A(SubCellInput2[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n19) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U1 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n26), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n25), .ZN(Red_MCInst2_MC0_v0_2[2]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U9 ( .A1(SubCellInput2[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n27), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n28) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U8 ( .A1(SubCellInput2[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n26), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n27) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_2_U7 ( .A(SubCellInput2[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n26) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n25), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n24), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n29) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U5 ( .A(
        SubCellInst2_LFInst_15_LFInst_2_n23), .B(SubCellInput2[62]), .Z(
        SubCellInst2_LFInst_15_LFInst_2_n24) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U4 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n23) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n22), .A2(SubCellInput2[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n25) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U2 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n22) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U1 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n29), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n28), .ZN(MCInst2_MC0_v0_3[3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U9 ( .A1(SubCellInput2[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n24), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n25) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U8 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n23), .A2(SubCellInput2[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n24) );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_3_U7 ( .A1(SubCellInput2[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n22), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n26) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n23), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n21), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n22) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U5 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n20), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n19), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n21) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U4 ( .A1(SubCellInput2[62]), .A2(
        SubCellInput2[60]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n19) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_3_U3 ( .A(SubCellInput2[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n20) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U2 ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n23) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U1 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n26), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n25), .ZN(Red_MCInst2_MC0_v0_1[0]) );
  BUF_X1 MCInst2_MC0_U2 ( .A(ShiftRowsOutput2[28]), .Z(MCInst2_MC0_v2_3[1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U2 ( .A(MCInst2_MC0_v0_2Inst_0_n3), .B(
        Red_MCInst2_MC0_v0_1[0]), .ZN(MCInst2_MC0_v0_2[0]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_2[2]), .ZN(MCInst2_MC0_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_0_U1 ( .A(MCInst2_MC0_v1_3[3]), .B(
        Red_MCInst2_MC0_v1_1[2]), .Z(MCInst2_MC0_v1_1[0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U2 ( .A(MCInst2_MC0_v1_2Inst_0_n3), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_v1_2[0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U1 ( .A(MCInst2_MC0_v1_3[2]), .B(
        MCInst2_MC0_v1_3[3]), .ZN(MCInst2_MC0_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_0_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[3]), .Z(MCInst2_MC0_v2_1[0]) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_0_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        Red_MCInst2_MC0_v2_2[1]), .Z(MCInst2_MC0_v2_2[0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U3 ( .A(MCInst2_MC0_v2_3Inst_0_n6), .B(
        MCInst2_MC0_v2_3Inst_0_n5), .ZN(MCInst2_MC0_v2_3[0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(MCInst2_MC0_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_0_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(MCInst2_MC0_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_0_U1 ( .A(MCInst2_MC0_v3_0[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_v3_1[0]) );
  XOR2_X1 MCInst2_MC0_v3_2Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(MCInst2_MC0_v3_2[0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U2 ( .A(MCInst2_MC0_v3_3Inst_0_n3), .B(
        Red_MCInst2_MC0_v3_1[2]), .ZN(MCInst2_MC0_v3_3[0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .ZN(MCInst2_MC0_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_1_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(MCInst2_MC0_v0_0[1]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), .B(
        MCInst2_MC0_v0_3[3]), .Z(MCInst2_MC0_v0_1[1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U2 ( .A(MCInst2_MC0_v0_2Inst_1_n3), .B(
        Red_MCInst2_MC0_v0_1[0]), .ZN(MCInst2_MC0_v0_2[1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        MCInst2_MC0_v0_3[3]), .ZN(MCInst2_MC0_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(MCInst2_MC0_v0_3[1]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        MCInst2_MC0_v1_3[3]), .Z(MCInst2_MC0_v1_1[1]) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        MCInst2_MC0_v1_3[2]), .Z(MCInst2_MC0_v1_2[1]) );
  XOR2_X1 MCInst2_MC0_v1_3Inst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_1[2]), .Z(MCInst2_MC0_v1_3[1]) );
  XOR2_X1 MCInst2_MC0_v2_0Inst_1_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        Red_MCInst2_MC0_v2_2[1]), .Z(MCInst2_MC0_v2_0[1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U2 ( .A(MCInst2_MC0_v2_1Inst_1_n3), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(MCInst2_MC0_v2_1[1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U3 ( .A(MCInst2_MC0_v2_2Inst_1_n6), .B(
        MCInst2_MC0_v2_2Inst_1_n5), .ZN(MCInst2_MC0_v2_2[1]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(MCInst2_MC0_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_1_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(MCInst2_MC0_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC0_v3_0Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_v3_0[1]) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[3]), .Z(MCInst2_MC0_v3_1[1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U2 ( .A(MCInst2_MC0_v3_3Inst_1_n3), .B(
        Red_MCInst2_MC0_v3_1[2]), .ZN(MCInst2_MC0_v3_3[1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[3]), .ZN(MCInst2_MC0_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(MCInst2_MC0_v0_0[2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_2_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(MCInst2_MC0_v0_1[2]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_2_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(MCInst2_MC0_v0_2[2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U2 ( .A(MCInst2_MC0_v1_1Inst_2_n3), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_v1_1[2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U2 ( .A(MCInst2_MC0_v1_2Inst_2_n3), .B(
        MCInst2_MC0_v1_3[3]), .ZN(MCInst2_MC0_v1_2[2]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U2 ( .A(MCInst2_MC0_v2_1Inst_2_n3), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(MCInst2_MC0_v2_1[2]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U2 ( .A(MCInst2_MC0_v2_2Inst_2_n3), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(MCInst2_MC0_v2_2[2]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_2_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(MCInst2_MC0_v2_3[2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U2 ( .A(MCInst2_MC0_v3_1Inst_2_n3), .B(
        Red_MCInst2_MC0_v3_1[2]), .ZN(MCInst2_MC0_v3_1[2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .ZN(MCInst2_MC0_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_2_U1 ( .A(Red_MCInst2_MC0_v3_3[2]), .B(
        Red_MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_v3_3[2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(MCInst2_MC0_v0_1[3]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        MCInst2_MC0_v0_3[3]), .Z(MCInst2_MC0_v0_2[3]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_3_U1 ( .A(MCInst2_MC0_v1_3[2]), .B(
        MCInst2_MC0_v1_3[3]), .Z(MCInst2_MC0_v1_1[3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U3 ( .A(MCInst2_MC0_v1_2Inst_3_n6), .B(
        MCInst2_MC0_v1_2Inst_3_n5), .ZN(MCInst2_MC0_v1_2[3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U2 ( .A(MCInst2_MC0_v1_3[3]), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_3_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        MCInst2_MC0_v1_3[2]), .Z(MCInst2_MC0_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_3_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        Red_MCInst2_MC0_v2_2[1]), .Z(MCInst2_MC0_v2_1[3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U2 ( .A(MCInst2_MC0_v2_2Inst_3_n3), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(MCInst2_MC0_v2_2[3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U2 ( .A(MCInst2_MC0_v2_3Inst_3_n3), .B(
        MCInst2_MC0_v2_0[3]), .ZN(MCInst2_MC0_v2_3[3]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U1 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v2_0[2]), .ZN(MCInst2_MC0_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_3_U1 ( .A(Red_MCInst2_MC0_v3_3[2]), .B(
        MCInst2_MC0_v3_0[3]), .Z(MCInst2_MC0_v3_1[3]) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_3_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[3]), .Z(MCInst2_MC0_v3_3[3]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[60]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_2[1]), 
        .B(MCInst2_MC0_v1_0_0_), .ZN(MCInst2_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[61]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_0[1]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_0[1]), .B(
        MCInst2_MC0_v3_0[1]), .Z(MCInst2_MC0_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[62]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v1_3[3]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_0[2]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(MCInst2_MC0_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[63]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), .B(
        MCInst2_MC0_v3_0[3]), .Z(MCInst2_MC0_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[44]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_1[0]), .B(
        MCInst2_MC0_v1_1[0]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), .B(
        MCInst2_MC0_v3_1[0]), .Z(MCInst2_MC0_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[45]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v1_1[1]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_1[1]), .B(
        MCInst2_MC0_v3_1[1]), .Z(MCInst2_MC0_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[46]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_1[2]), .B(
        MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_1[2]), .B(
        MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[47]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_1[3]), .B(
        MCInst2_MC0_v1_1[3]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_1[3]), .B(
        MCInst2_MC0_v3_1[3]), .Z(MCInst2_MC0_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[28]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_2[0]), .B(
        MCInst2_MC0_v1_2[0]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC0_v0_2[0]), .B(
        MCInst2_MC0_v3_2[0]), .Z(MCInst2_MC0_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[29]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_2[1]), .B(
        MCInst2_MC0_v1_2[1]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_2[1]), .B(
        MCInst2_MC0_v3_0[3]), .Z(MCInst2_MC0_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[30]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_2[2]), .B(
        MCInst2_MC0_v1_2[2]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC0_v0_2[2]), .B(
        Red_MCInst2_MC0_v3_1[2]), .Z(MCInst2_MC0_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[31]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_2[3]), .B(
        MCInst2_MC0_v1_2[3]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_2[3]), .B(
        MCInst2_MC0_v3_2[3]), .Z(MCInst2_MC0_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[12]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC0_v2_3[0]), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_1[0]), .B(
        MCInst2_MC0_v3_3[0]), .Z(MCInst2_MC0_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[13]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC0_v2_3[1]), .B(
        MCInst2_MC0_v1_3[1]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC0_v0_3[1]), .B(
        MCInst2_MC0_v3_3[1]), .Z(MCInst2_MC0_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[14]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC0_v2_3[2]), .B(
        MCInst2_MC0_v1_3[2]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), .B(
        MCInst2_MC0_v3_3[2]), .Z(MCInst2_MC0_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC0_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[15]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC0_v2_3[3]), .B(
        MCInst2_MC0_v1_3[3]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        MCInst2_MC0_v3_3[3]), .Z(MCInst2_MC0_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst2_MC1_U2 ( .A(ShiftRowsOutput2[24]), .Z(MCInst2_MC1_v2_3[1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U2 ( .A(MCInst2_MC1_v0_2Inst_0_n3), .B(
        Red_MCInst2_MC1_v0_1[0]), .ZN(MCInst2_MC1_v0_2[0]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_2[2]), .ZN(MCInst2_MC1_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_0_U1 ( .A(MCInst2_MC1_v1_3[3]), .B(
        Red_MCInst2_MC1_v1_1[2]), .Z(MCInst2_MC1_v1_1[0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U2 ( .A(MCInst2_MC1_v1_2Inst_0_n3), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_v1_2[0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U1 ( .A(MCInst2_MC1_v1_3[2]), .B(
        MCInst2_MC1_v1_3[3]), .ZN(MCInst2_MC1_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_0_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[3]), .Z(MCInst2_MC1_v2_1[0]) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_0_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        Red_MCInst2_MC1_v2_2[1]), .Z(MCInst2_MC1_v2_2[0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U3 ( .A(MCInst2_MC1_v2_3Inst_0_n6), .B(
        MCInst2_MC1_v2_3Inst_0_n5), .ZN(MCInst2_MC1_v2_3[0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(MCInst2_MC1_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_0_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(MCInst2_MC1_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_0_U1 ( .A(MCInst2_MC1_v3_0[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_v3_1[0]) );
  XOR2_X1 MCInst2_MC1_v3_2Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(MCInst2_MC1_v3_2[0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U2 ( .A(MCInst2_MC1_v3_3Inst_0_n3), .B(
        Red_MCInst2_MC1_v3_1[2]), .ZN(MCInst2_MC1_v3_3[0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .ZN(MCInst2_MC1_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_1_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(MCInst2_MC1_v0_0[1]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), .B(
        MCInst2_MC1_v0_3[3]), .Z(MCInst2_MC1_v0_1[1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U2 ( .A(MCInst2_MC1_v0_2Inst_1_n3), .B(
        Red_MCInst2_MC1_v0_1[0]), .ZN(MCInst2_MC1_v0_2[1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        MCInst2_MC1_v0_3[3]), .ZN(MCInst2_MC1_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(MCInst2_MC1_v0_3[1]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        MCInst2_MC1_v1_3[3]), .Z(MCInst2_MC1_v1_1[1]) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        MCInst2_MC1_v1_3[2]), .Z(MCInst2_MC1_v1_2[1]) );
  XOR2_X1 MCInst2_MC1_v1_3Inst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_1[2]), .Z(MCInst2_MC1_v1_3[1]) );
  XOR2_X1 MCInst2_MC1_v2_0Inst_1_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        Red_MCInst2_MC1_v2_2[1]), .Z(MCInst2_MC1_v2_0[1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U2 ( .A(MCInst2_MC1_v2_1Inst_1_n3), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(MCInst2_MC1_v2_1[1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U3 ( .A(MCInst2_MC1_v2_2Inst_1_n6), .B(
        MCInst2_MC1_v2_2Inst_1_n5), .ZN(MCInst2_MC1_v2_2[1]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(MCInst2_MC1_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_1_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(MCInst2_MC1_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC1_v3_0Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_v3_0[1]) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[3]), .Z(MCInst2_MC1_v3_1[1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U2 ( .A(MCInst2_MC1_v3_3Inst_1_n3), .B(
        Red_MCInst2_MC1_v3_1[2]), .ZN(MCInst2_MC1_v3_3[1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[3]), .ZN(MCInst2_MC1_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(MCInst2_MC1_v0_0[2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_2_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(MCInst2_MC1_v0_1[2]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_2_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(MCInst2_MC1_v0_2[2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U2 ( .A(MCInst2_MC1_v1_1Inst_2_n3), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_v1_1[2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U2 ( .A(MCInst2_MC1_v1_2Inst_2_n3), .B(
        MCInst2_MC1_v1_3[3]), .ZN(MCInst2_MC1_v1_2[2]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U2 ( .A(MCInst2_MC1_v2_1Inst_2_n3), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(MCInst2_MC1_v2_1[2]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U2 ( .A(MCInst2_MC1_v2_2Inst_2_n3), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(MCInst2_MC1_v2_2[2]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_2_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(MCInst2_MC1_v2_3[2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U2 ( .A(MCInst2_MC1_v3_1Inst_2_n3), .B(
        Red_MCInst2_MC1_v3_1[2]), .ZN(MCInst2_MC1_v3_1[2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .ZN(MCInst2_MC1_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_2_U1 ( .A(Red_MCInst2_MC1_v3_3[2]), .B(
        Red_MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_v3_3[2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(MCInst2_MC1_v0_1[3]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        MCInst2_MC1_v0_3[3]), .Z(MCInst2_MC1_v0_2[3]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_3_U1 ( .A(MCInst2_MC1_v1_3[2]), .B(
        MCInst2_MC1_v1_3[3]), .Z(MCInst2_MC1_v1_1[3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U3 ( .A(MCInst2_MC1_v1_2Inst_3_n6), .B(
        MCInst2_MC1_v1_2Inst_3_n5), .ZN(MCInst2_MC1_v1_2[3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U2 ( .A(MCInst2_MC1_v1_3[3]), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_3_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        MCInst2_MC1_v1_3[2]), .Z(MCInst2_MC1_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_3_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        Red_MCInst2_MC1_v2_2[1]), .Z(MCInst2_MC1_v2_1[3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U2 ( .A(MCInst2_MC1_v2_2Inst_3_n3), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(MCInst2_MC1_v2_2[3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U2 ( .A(MCInst2_MC1_v2_3Inst_3_n3), .B(
        MCInst2_MC1_v2_0[3]), .ZN(MCInst2_MC1_v2_3[3]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U1 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v2_0[2]), .ZN(MCInst2_MC1_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_3_U1 ( .A(Red_MCInst2_MC1_v3_3[2]), .B(
        MCInst2_MC1_v3_0[3]), .Z(MCInst2_MC1_v3_1[3]) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_3_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[3]), .Z(MCInst2_MC1_v3_3[3]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[56]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_2[1]), 
        .B(MCInst2_MC1_v1_0_0_), .ZN(MCInst2_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[57]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_0[1]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_0[1]), .B(
        MCInst2_MC1_v3_0[1]), .Z(MCInst2_MC1_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[58]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v1_3[3]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_0[2]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(MCInst2_MC1_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[59]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), .B(
        MCInst2_MC1_v3_0[3]), .Z(MCInst2_MC1_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[40]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_1[0]), .B(
        MCInst2_MC1_v1_1[0]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), .B(
        MCInst2_MC1_v3_1[0]), .Z(MCInst2_MC1_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[41]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v1_1[1]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_1[1]), .B(
        MCInst2_MC1_v3_1[1]), .Z(MCInst2_MC1_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[42]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_1[2]), .B(
        MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_1[2]), .B(
        MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[43]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_1[3]), .B(
        MCInst2_MC1_v1_1[3]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_1[3]), .B(
        MCInst2_MC1_v3_1[3]), .Z(MCInst2_MC1_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[24]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_2[0]), .B(
        MCInst2_MC1_v1_2[0]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC1_v0_2[0]), .B(
        MCInst2_MC1_v3_2[0]), .Z(MCInst2_MC1_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[25]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_2[1]), .B(
        MCInst2_MC1_v1_2[1]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_2[1]), .B(
        MCInst2_MC1_v3_0[3]), .Z(MCInst2_MC1_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[26]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_2[2]), .B(
        MCInst2_MC1_v1_2[2]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC1_v0_2[2]), .B(
        Red_MCInst2_MC1_v3_1[2]), .Z(MCInst2_MC1_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[27]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_2[3]), .B(
        MCInst2_MC1_v1_2[3]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_2[3]), .B(
        MCInst2_MC1_v3_2[3]), .Z(MCInst2_MC1_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[8]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC1_v2_3[0]), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_1[0]), .B(
        MCInst2_MC1_v3_3[0]), .Z(MCInst2_MC1_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[9]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC1_v2_3[1]), .B(
        MCInst2_MC1_v1_3[1]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC1_v0_3[1]), .B(
        MCInst2_MC1_v3_3[1]), .Z(MCInst2_MC1_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[10]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC1_v2_3[2]), .B(
        MCInst2_MC1_v1_3[2]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), .B(
        MCInst2_MC1_v3_3[2]), .Z(MCInst2_MC1_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC1_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[11]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC1_v2_3[3]), .B(
        MCInst2_MC1_v1_3[3]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        MCInst2_MC1_v3_3[3]), .Z(MCInst2_MC1_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst2_MC2_U2 ( .A(ShiftRowsOutput2[20]), .Z(MCInst2_MC2_v2_3[1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U2 ( .A(MCInst2_MC2_v0_2Inst_0_n3), .B(
        Red_MCInst2_MC2_v0_1[0]), .ZN(MCInst2_MC2_v0_2[0]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_2[2]), .ZN(MCInst2_MC2_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_0_U1 ( .A(MCInst2_MC2_v1_3[3]), .B(
        Red_MCInst2_MC2_v1_1[2]), .Z(MCInst2_MC2_v1_1[0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U2 ( .A(MCInst2_MC2_v1_2Inst_0_n3), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_v1_2[0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U1 ( .A(MCInst2_MC2_v1_3[2]), .B(
        MCInst2_MC2_v1_3[3]), .ZN(MCInst2_MC2_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_0_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[3]), .Z(MCInst2_MC2_v2_1[0]) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_0_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        Red_MCInst2_MC2_v2_2[1]), .Z(MCInst2_MC2_v2_2[0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U3 ( .A(MCInst2_MC2_v2_3Inst_0_n6), .B(
        MCInst2_MC2_v2_3Inst_0_n5), .ZN(MCInst2_MC2_v2_3[0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(MCInst2_MC2_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_0_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(MCInst2_MC2_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_0_U1 ( .A(MCInst2_MC2_v3_0[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_v3_1[0]) );
  XOR2_X1 MCInst2_MC2_v3_2Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(MCInst2_MC2_v3_2[0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U2 ( .A(MCInst2_MC2_v3_3Inst_0_n3), .B(
        Red_MCInst2_MC2_v3_1[2]), .ZN(MCInst2_MC2_v3_3[0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .ZN(MCInst2_MC2_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_1_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(MCInst2_MC2_v0_0[1]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), .B(
        MCInst2_MC2_v0_3[3]), .Z(MCInst2_MC2_v0_1[1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U2 ( .A(MCInst2_MC2_v0_2Inst_1_n3), .B(
        Red_MCInst2_MC2_v0_1[0]), .ZN(MCInst2_MC2_v0_2[1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        MCInst2_MC2_v0_3[3]), .ZN(MCInst2_MC2_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(MCInst2_MC2_v0_3[1]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        MCInst2_MC2_v1_3[3]), .Z(MCInst2_MC2_v1_1[1]) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        MCInst2_MC2_v1_3[2]), .Z(MCInst2_MC2_v1_2[1]) );
  XOR2_X1 MCInst2_MC2_v1_3Inst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_1[2]), .Z(MCInst2_MC2_v1_3[1]) );
  XOR2_X1 MCInst2_MC2_v2_0Inst_1_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        Red_MCInst2_MC2_v2_2[1]), .Z(MCInst2_MC2_v2_0[1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U2 ( .A(MCInst2_MC2_v2_1Inst_1_n3), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(MCInst2_MC2_v2_1[1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U3 ( .A(MCInst2_MC2_v2_2Inst_1_n6), .B(
        MCInst2_MC2_v2_2Inst_1_n5), .ZN(MCInst2_MC2_v2_2[1]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(MCInst2_MC2_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_1_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(MCInst2_MC2_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC2_v3_0Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_v3_0[1]) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[3]), .Z(MCInst2_MC2_v3_1[1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U2 ( .A(MCInst2_MC2_v3_3Inst_1_n3), .B(
        Red_MCInst2_MC2_v3_1[2]), .ZN(MCInst2_MC2_v3_3[1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[3]), .ZN(MCInst2_MC2_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(MCInst2_MC2_v0_0[2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_2_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(MCInst2_MC2_v0_1[2]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_2_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(MCInst2_MC2_v0_2[2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U2 ( .A(MCInst2_MC2_v1_1Inst_2_n3), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_v1_1[2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U2 ( .A(MCInst2_MC2_v1_2Inst_2_n3), .B(
        MCInst2_MC2_v1_3[3]), .ZN(MCInst2_MC2_v1_2[2]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U2 ( .A(MCInst2_MC2_v2_1Inst_2_n3), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(MCInst2_MC2_v2_1[2]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U2 ( .A(MCInst2_MC2_v2_2Inst_2_n3), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(MCInst2_MC2_v2_2[2]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_2_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(MCInst2_MC2_v2_3[2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U2 ( .A(MCInst2_MC2_v3_1Inst_2_n3), .B(
        Red_MCInst2_MC2_v3_1[2]), .ZN(MCInst2_MC2_v3_1[2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .ZN(MCInst2_MC2_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_2_U1 ( .A(Red_MCInst2_MC2_v3_3[2]), .B(
        Red_MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_v3_3[2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(MCInst2_MC2_v0_1[3]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        MCInst2_MC2_v0_3[3]), .Z(MCInst2_MC2_v0_2[3]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_3_U1 ( .A(MCInst2_MC2_v1_3[2]), .B(
        MCInst2_MC2_v1_3[3]), .Z(MCInst2_MC2_v1_1[3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U3 ( .A(MCInst2_MC2_v1_2Inst_3_n6), .B(
        MCInst2_MC2_v1_2Inst_3_n5), .ZN(MCInst2_MC2_v1_2[3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U2 ( .A(MCInst2_MC2_v1_3[3]), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_3_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        MCInst2_MC2_v1_3[2]), .Z(MCInst2_MC2_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_3_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        Red_MCInst2_MC2_v2_2[1]), .Z(MCInst2_MC2_v2_1[3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U2 ( .A(MCInst2_MC2_v2_2Inst_3_n3), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(MCInst2_MC2_v2_2[3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U2 ( .A(MCInst2_MC2_v2_3Inst_3_n3), .B(
        MCInst2_MC2_v2_0[3]), .ZN(MCInst2_MC2_v2_3[3]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U1 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v2_0[2]), .ZN(MCInst2_MC2_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_3_U1 ( .A(Red_MCInst2_MC2_v3_3[2]), .B(
        MCInst2_MC2_v3_0[3]), .Z(MCInst2_MC2_v3_1[3]) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_3_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[3]), .Z(MCInst2_MC2_v3_3[3]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[52]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_2[1]), 
        .B(MCInst2_MC2_v1_0_0_), .ZN(MCInst2_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[53]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_0[1]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_0[1]), .B(
        MCInst2_MC2_v3_0[1]), .Z(MCInst2_MC2_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[54]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v1_3[3]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_0[2]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(MCInst2_MC2_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[55]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), .B(
        MCInst2_MC2_v3_0[3]), .Z(MCInst2_MC2_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[36]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_1[0]), .B(
        MCInst2_MC2_v1_1[0]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), .B(
        MCInst2_MC2_v3_1[0]), .Z(MCInst2_MC2_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[37]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v1_1[1]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_1[1]), .B(
        MCInst2_MC2_v3_1[1]), .Z(MCInst2_MC2_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[38]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_1[2]), .B(
        MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_1[2]), .B(
        MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[39]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_1[3]), .B(
        MCInst2_MC2_v1_1[3]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_1[3]), .B(
        MCInst2_MC2_v3_1[3]), .Z(MCInst2_MC2_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[20]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_2[0]), .B(
        MCInst2_MC2_v1_2[0]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC2_v0_2[0]), .B(
        MCInst2_MC2_v3_2[0]), .Z(MCInst2_MC2_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[21]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_2[1]), .B(
        MCInst2_MC2_v1_2[1]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_2[1]), .B(
        MCInst2_MC2_v3_0[3]), .Z(MCInst2_MC2_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[22]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_2[2]), .B(
        MCInst2_MC2_v1_2[2]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC2_v0_2[2]), .B(
        Red_MCInst2_MC2_v3_1[2]), .Z(MCInst2_MC2_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[23]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_2[3]), .B(
        MCInst2_MC2_v1_2[3]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_2[3]), .B(
        MCInst2_MC2_v3_2[3]), .Z(MCInst2_MC2_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[4]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC2_v2_3[0]), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_1[0]), .B(
        MCInst2_MC2_v3_3[0]), .Z(MCInst2_MC2_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[5]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC2_v2_3[1]), .B(
        MCInst2_MC2_v1_3[1]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC2_v0_3[1]), .B(
        MCInst2_MC2_v3_3[1]), .Z(MCInst2_MC2_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[6]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC2_v2_3[2]), .B(
        MCInst2_MC2_v1_3[2]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), .B(
        MCInst2_MC2_v3_3[2]), .Z(MCInst2_MC2_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC2_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[7]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC2_v2_3[3]), .B(
        MCInst2_MC2_v1_3[3]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        MCInst2_MC2_v3_3[3]), .Z(MCInst2_MC2_r3Inst_XORInst_0_3_n8) );
  BUF_X1 MCInst2_MC3_U2 ( .A(ShiftRowsOutput2[16]), .Z(MCInst2_MC3_v2_3[1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U2 ( .A(MCInst2_MC3_v0_2Inst_0_n3), .B(
        Red_MCInst2_MC3_v0_1[0]), .ZN(MCInst2_MC3_v0_2[0]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_2[2]), .ZN(MCInst2_MC3_v0_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_0_U1 ( .A(MCInst2_MC3_v1_3[3]), .B(
        Red_MCInst2_MC3_v1_1[2]), .Z(MCInst2_MC3_v1_1[0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U2 ( .A(MCInst2_MC3_v1_2Inst_0_n3), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_v1_2[0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U1 ( .A(MCInst2_MC3_v1_3[2]), .B(
        MCInst2_MC3_v1_3[3]), .ZN(MCInst2_MC3_v1_2Inst_0_n3) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_0_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[3]), .Z(MCInst2_MC3_v2_1[0]) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_0_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        Red_MCInst2_MC3_v2_2[1]), .Z(MCInst2_MC3_v2_2[0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U3 ( .A(MCInst2_MC3_v2_3Inst_0_n6), .B(
        MCInst2_MC3_v2_3Inst_0_n5), .ZN(MCInst2_MC3_v2_3[0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(MCInst2_MC3_v2_3Inst_0_n5) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_0_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(MCInst2_MC3_v2_3Inst_0_n6) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_0_U1 ( .A(MCInst2_MC3_v3_0[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_v3_1[0]) );
  XOR2_X1 MCInst2_MC3_v3_2Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(MCInst2_MC3_v3_2[0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U2 ( .A(MCInst2_MC3_v3_3Inst_0_n3), .B(
        Red_MCInst2_MC3_v3_1[2]), .ZN(MCInst2_MC3_v3_3[0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .ZN(MCInst2_MC3_v3_3Inst_0_n3) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_1_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(MCInst2_MC3_v0_0[1]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), .B(
        MCInst2_MC3_v0_3[3]), .Z(MCInst2_MC3_v0_1[1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U2 ( .A(MCInst2_MC3_v0_2Inst_1_n3), .B(
        Red_MCInst2_MC3_v0_1[0]), .ZN(MCInst2_MC3_v0_2[1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        MCInst2_MC3_v0_3[3]), .ZN(MCInst2_MC3_v0_2Inst_1_n3) );
  XOR2_X1 MCInst2_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(MCInst2_MC3_v0_3[1]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        MCInst2_MC3_v1_3[3]), .Z(MCInst2_MC3_v1_1[1]) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        MCInst2_MC3_v1_3[2]), .Z(MCInst2_MC3_v1_2[1]) );
  XOR2_X1 MCInst2_MC3_v1_3Inst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_1[2]), .Z(MCInst2_MC3_v1_3[1]) );
  XOR2_X1 MCInst2_MC3_v2_0Inst_1_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        Red_MCInst2_MC3_v2_2[1]), .Z(MCInst2_MC3_v2_0[1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U2 ( .A(MCInst2_MC3_v2_1Inst_1_n3), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(MCInst2_MC3_v2_1[1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_1Inst_1_n3) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U3 ( .A(MCInst2_MC3_v2_2Inst_1_n6), .B(
        MCInst2_MC3_v2_2Inst_1_n5), .ZN(MCInst2_MC3_v2_2[1]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(MCInst2_MC3_v2_2Inst_1_n5) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_1_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(MCInst2_MC3_v2_2Inst_1_n6) );
  XOR2_X1 MCInst2_MC3_v3_0Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_v3_0[1]) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[3]), .Z(MCInst2_MC3_v3_1[1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U2 ( .A(MCInst2_MC3_v3_3Inst_1_n3), .B(
        Red_MCInst2_MC3_v3_1[2]), .ZN(MCInst2_MC3_v3_3[1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[3]), .ZN(MCInst2_MC3_v3_3Inst_1_n3) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(MCInst2_MC3_v0_0[2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_2_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(MCInst2_MC3_v0_1[2]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_2_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(MCInst2_MC3_v0_2[2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U2 ( .A(MCInst2_MC3_v1_1Inst_2_n3), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_v1_1[2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_v1_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U2 ( .A(MCInst2_MC3_v1_2Inst_2_n3), .B(
        MCInst2_MC3_v1_3[3]), .ZN(MCInst2_MC3_v1_2[2]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U2 ( .A(MCInst2_MC3_v2_1Inst_2_n3), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(MCInst2_MC3_v2_1[2]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_1Inst_2_n3) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U2 ( .A(MCInst2_MC3_v2_2Inst_2_n3), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(MCInst2_MC3_v2_2[2]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_2Inst_2_n3) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_2_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(MCInst2_MC3_v2_3[2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U2 ( .A(MCInst2_MC3_v3_1Inst_2_n3), .B(
        Red_MCInst2_MC3_v3_1[2]), .ZN(MCInst2_MC3_v3_1[2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .ZN(MCInst2_MC3_v3_1Inst_2_n3) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_2_U1 ( .A(Red_MCInst2_MC3_v3_3[2]), .B(
        Red_MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_v3_3[2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_3_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(MCInst2_MC3_v0_1[3]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_3_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        MCInst2_MC3_v0_3[3]), .Z(MCInst2_MC3_v0_2[3]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_3_U1 ( .A(MCInst2_MC3_v1_3[2]), .B(
        MCInst2_MC3_v1_3[3]), .Z(MCInst2_MC3_v1_1[3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U3 ( .A(MCInst2_MC3_v1_2Inst_3_n6), .B(
        MCInst2_MC3_v1_2Inst_3_n5), .ZN(MCInst2_MC3_v1_2[3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U2 ( .A(MCInst2_MC3_v1_3[3]), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_v1_2Inst_3_n5) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_3_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        MCInst2_MC3_v1_3[2]), .Z(MCInst2_MC3_v1_2Inst_3_n6) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_3_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        Red_MCInst2_MC3_v2_2[1]), .Z(MCInst2_MC3_v2_1[3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U2 ( .A(MCInst2_MC3_v2_2Inst_3_n3), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(MCInst2_MC3_v2_2[3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_2Inst_3_n3) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U2 ( .A(MCInst2_MC3_v2_3Inst_3_n3), .B(
        MCInst2_MC3_v2_0[3]), .ZN(MCInst2_MC3_v2_3[3]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U1 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v2_0[2]), .ZN(MCInst2_MC3_v2_3Inst_3_n3) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_3_U1 ( .A(Red_MCInst2_MC3_v3_3[2]), .B(
        MCInst2_MC3_v3_0[3]), .Z(MCInst2_MC3_v3_1[3]) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_3_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[3]), .Z(MCInst2_MC3_v3_3[3]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_0_n7), .ZN(Ciphertext[48]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_2[1]), 
        .B(MCInst2_MC3_v1_0_0_), .ZN(MCInst2_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_r0Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_1_n7), .ZN(Ciphertext[49]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_0[1]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_0[1]), .B(
        MCInst2_MC3_v3_0[1]), .Z(MCInst2_MC3_r0Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_2_n7), .ZN(Ciphertext[50]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v1_3[3]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_0[2]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(MCInst2_MC3_r0Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r0Inst_XORInst_0_3_n7), .ZN(Ciphertext[51]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), .B(
        MCInst2_MC3_v3_0[3]), .Z(MCInst2_MC3_r0Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_0_n7), .ZN(Ciphertext[32]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_1[0]), .B(
        MCInst2_MC3_v1_1[0]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), .B(
        MCInst2_MC3_v3_1[0]), .Z(MCInst2_MC3_r1Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_1_n7), .ZN(Ciphertext[33]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v1_1[1]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_1[1]), .B(
        MCInst2_MC3_v3_1[1]), .Z(MCInst2_MC3_r1Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_2_n7), .ZN(Ciphertext[34]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_1[2]), .B(
        MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_1[2]), .B(
        MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_r1Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r1Inst_XORInst_0_3_n7), .ZN(Ciphertext[35]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_1[3]), .B(
        MCInst2_MC3_v1_1[3]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_1[3]), .B(
        MCInst2_MC3_v3_1[3]), .Z(MCInst2_MC3_r1Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_0_n7), .ZN(Ciphertext[16]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_2[0]), .B(
        MCInst2_MC3_v1_2[0]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U1 ( .A(MCInst2_MC3_v0_2[0]), .B(
        MCInst2_MC3_v3_2[0]), .Z(MCInst2_MC3_r2Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_1_n7), .ZN(Ciphertext[17]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_2[1]), .B(
        MCInst2_MC3_v1_2[1]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_2[1]), .B(
        MCInst2_MC3_v3_0[3]), .Z(MCInst2_MC3_r2Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_2_n7), .ZN(Ciphertext[18]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_2[2]), .B(
        MCInst2_MC3_v1_2[2]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U1 ( .A(MCInst2_MC3_v0_2[2]), .B(
        Red_MCInst2_MC3_v3_1[2]), .Z(MCInst2_MC3_r2Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r2Inst_XORInst_0_3_n7), .ZN(Ciphertext[19]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_2[3]), .B(
        MCInst2_MC3_v1_2[3]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_2[3]), .B(
        MCInst2_MC3_v3_2[3]), .Z(MCInst2_MC3_r2Inst_XORInst_0_3_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_0_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_0_n7), .ZN(Ciphertext[0]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U2 ( .A(MCInst2_MC3_v2_3[0]), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_1[0]), .B(
        MCInst2_MC3_v3_3[0]), .Z(MCInst2_MC3_r3Inst_XORInst_0_0_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_1_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_1_n7), .ZN(Ciphertext[1]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U2 ( .A(MCInst2_MC3_v2_3[1]), .B(
        MCInst2_MC3_v1_3[1]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U1 ( .A(MCInst2_MC3_v0_3[1]), .B(
        MCInst2_MC3_v3_3[1]), .Z(MCInst2_MC3_r3Inst_XORInst_0_1_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_2_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_2_n7), .ZN(Ciphertext[2]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U2 ( .A(MCInst2_MC3_v2_3[2]), .B(
        MCInst2_MC3_v1_3[2]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), .B(
        MCInst2_MC3_v3_3[2]), .Z(MCInst2_MC3_r3Inst_XORInst_0_2_n8) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U3 ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_3_n8), .B(
        MCInst2_MC3_r3Inst_XORInst_0_3_n7), .ZN(Ciphertext[3]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U2 ( .A(MCInst2_MC3_v2_3[3]), .B(
        MCInst2_MC3_v1_3[3]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_3_n7) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        MCInst2_MC3_v3_3[3]), .Z(MCInst2_MC3_r3Inst_XORInst_0_3_n8) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n3), .B(Plaintext[2]), .ZN(
        Red_Plaintext[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Plaintext[0]), .B(
        Plaintext[1]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_1_n3), .B(Plaintext[3]), .ZN(
        Red_Plaintext[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U1 ( .A(Plaintext[0]), .B(
        Plaintext[1]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_2_n3), .B(Plaintext[3]), .ZN(
        Red_Plaintext[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U1 ( .A(Plaintext[1]), .B(
        Plaintext[2]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n3), .B(Plaintext[6]), .ZN(
        Red_Plaintext[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Plaintext[4]), .B(
        Plaintext[5]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_1_n3), .B(Plaintext[7]), .ZN(
        Red_Plaintext[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U1 ( .A(Plaintext[4]), .B(
        Plaintext[5]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_2_n3), .B(Plaintext[7]), .ZN(
        Red_Plaintext[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U1 ( .A(Plaintext[5]), .B(
        Plaintext[6]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n3), .B(Plaintext[10]), .ZN(
        Red_Plaintext[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Plaintext[8]), .B(
        Plaintext[9]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_1_n3), .B(Plaintext[11]), .ZN(
        Red_Plaintext[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U1 ( .A(Plaintext[8]), .B(
        Plaintext[9]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_2_n3), .B(Plaintext[11]), .ZN(
        Red_Plaintext[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U1 ( .A(Plaintext[9]), .B(
        Plaintext[10]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n3), .B(Plaintext[14]), .ZN(
        Red_Plaintext[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Plaintext[12]), .B(
        Plaintext[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_1_n3), .B(Plaintext[15]), .ZN(
        Red_Plaintext[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U1 ( .A(Plaintext[12]), .B(
        Plaintext[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_2_n3), .B(Plaintext[15]), .ZN(
        Red_Plaintext[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U1 ( .A(Plaintext[13]), .B(
        Plaintext[14]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n3), .B(Plaintext[18]), .ZN(
        Red_Plaintext[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Plaintext[16]), .B(
        Plaintext[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_1_n3), .B(Plaintext[19]), .ZN(
        Red_Plaintext[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U1 ( .A(Plaintext[16]), .B(
        Plaintext[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_2_n3), .B(Plaintext[19]), .ZN(
        Red_Plaintext[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U1 ( .A(Plaintext[17]), .B(
        Plaintext[18]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n3), .B(Plaintext[22]), .ZN(
        Red_Plaintext[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Plaintext[20]), .B(
        Plaintext[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_1_n3), .B(Plaintext[23]), .ZN(
        Red_Plaintext[16]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U1 ( .A(Plaintext[20]), .B(
        Plaintext[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_2_n3), .B(Plaintext[23]), .ZN(
        Red_Plaintext[17]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U1 ( .A(Plaintext[21]), .B(
        Plaintext[22]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n3), .B(Plaintext[26]), .ZN(
        Red_Plaintext[18]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Plaintext[24]), .B(
        Plaintext[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_1_n3), .B(Plaintext[27]), .ZN(
        Red_Plaintext[19]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U1 ( .A(Plaintext[24]), .B(
        Plaintext[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_2_n3), .B(Plaintext[27]), .ZN(
        Red_Plaintext[20]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U1 ( .A(Plaintext[25]), .B(
        Plaintext[26]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n3), .B(Plaintext[30]), .ZN(
        Red_Plaintext[21]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Plaintext[28]), .B(
        Plaintext[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_1_n3), .B(Plaintext[31]), .ZN(
        Red_Plaintext[22]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U1 ( .A(Plaintext[28]), .B(
        Plaintext[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_2_n3), .B(Plaintext[31]), .ZN(
        Red_Plaintext[23]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U1 ( .A(Plaintext[29]), .B(
        Plaintext[30]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n3), .B(Plaintext[34]), .ZN(
        Red_Plaintext[24]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Plaintext[32]), .B(
        Plaintext[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_1_n3), .B(Plaintext[35]), .ZN(
        Red_Plaintext[25]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U1 ( .A(Plaintext[32]), .B(
        Plaintext[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_2_n3), .B(Plaintext[35]), .ZN(
        Red_Plaintext[26]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U1 ( .A(Plaintext[33]), .B(
        Plaintext[34]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n3), .B(Plaintext[38]), .ZN(
        Red_Plaintext[27]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Plaintext[36]), .B(
        Plaintext[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_1_n3), .B(Plaintext[39]), .ZN(
        Red_Plaintext[28]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U1 ( .A(Plaintext[36]), .B(
        Plaintext[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_2_n3), .B(Plaintext[39]), .ZN(
        Red_Plaintext[29]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U1 ( .A(Plaintext[37]), .B(
        Plaintext[38]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n3), .B(Plaintext[42]), .ZN(
        Red_Plaintext[30]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Plaintext[40]), .B(
        Plaintext[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_1_n3), .B(Plaintext[43]), .ZN(
        Red_Plaintext[31]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U1 ( .A(Plaintext[40]), .B(
        Plaintext[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_2_n3), .B(Plaintext[43]), .ZN(
        Red_Plaintext[32]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U1 ( .A(Plaintext[41]), .B(
        Plaintext[42]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n3), .B(Plaintext[46]), .ZN(
        Red_Plaintext[33]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Plaintext[44]), .B(
        Plaintext[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_1_n3), .B(Plaintext[47]), .ZN(
        Red_Plaintext[34]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U1 ( .A(Plaintext[44]), .B(
        Plaintext[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_2_n3), .B(Plaintext[47]), .ZN(
        Red_Plaintext[35]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U1 ( .A(Plaintext[45]), .B(
        Plaintext[46]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n3), .B(Plaintext[50]), .ZN(
        Red_Plaintext[36]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Plaintext[48]), .B(
        Plaintext[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_1_n3), .B(Plaintext[51]), .ZN(
        Red_Plaintext[37]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U1 ( .A(Plaintext[48]), .B(
        Plaintext[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_2_n3), .B(Plaintext[51]), .ZN(
        Red_Plaintext[38]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U1 ( .A(Plaintext[49]), .B(
        Plaintext[50]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n3), .B(Plaintext[54]), .ZN(
        Red_Plaintext[39]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Plaintext[52]), .B(
        Plaintext[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_1_n3), .B(Plaintext[55]), .ZN(
        Red_Plaintext[40]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U1 ( .A(Plaintext[52]), .B(
        Plaintext[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_2_n3), .B(Plaintext[55]), .ZN(
        Red_Plaintext[41]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U1 ( .A(Plaintext[53]), .B(
        Plaintext[54]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n3), .B(Plaintext[58]), .ZN(
        Red_Plaintext[42]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Plaintext[56]), .B(
        Plaintext[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_1_n3), .B(Plaintext[59]), .ZN(
        Red_Plaintext[43]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U1 ( .A(Plaintext[56]), .B(
        Plaintext[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_2_n3), .B(Plaintext[59]), .ZN(
        Red_Plaintext[44]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U1 ( .A(Plaintext[57]), .B(
        Plaintext[58]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n3), .B(Plaintext[62]), .ZN(
        Red_Plaintext[45]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Plaintext[60]), .B(
        Plaintext[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_1_n3), .B(Plaintext[63]), .ZN(
        Red_Plaintext[46]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U1 ( .A(Plaintext[60]), .B(
        Plaintext[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_2_n3), .B(Plaintext[63]), .ZN(
        Red_Plaintext[47]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U1 ( .A(Plaintext[61]), .B(
        Plaintext[62]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_2_n3) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_0_U1 ( .A(Red_Plaintext[0]), .B(
        Red_RoundKey[0]), .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_1_U1 ( .A(Red_Plaintext[1]), .B(
        Red_RoundKey[1]), .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_2_U1 ( .A(Red_Plaintext[2]), .B(
        Red_RoundKey[2]), .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_0_U1 ( .A(Red_Plaintext[3]), .B(
        Red_RoundKey[3]), .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_1_U1 ( .A(Red_Plaintext[4]), .B(
        Red_RoundKey[4]), .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_2_U1 ( .A(Red_Plaintext[5]), .B(
        Red_RoundKey[5]), .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_0_U1 ( .A(Red_Plaintext[6]), .B(
        Red_RoundKey[6]), .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_1_U1 ( .A(Red_Plaintext[7]), .B(
        Red_RoundKey[7]), .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_2_U1 ( .A(Red_Plaintext[8]), .B(
        Red_RoundKey[8]), .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_0_U1 ( .A(Red_Plaintext[9]), .B(
        Red_RoundKey[9]), .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_1_U1 ( .A(Red_Plaintext[10]), .B(
        Red_RoundKey[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_2_U1 ( .A(Red_Plaintext[11]), .B(
        Red_RoundKey[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_0_U1 ( .A(Red_Plaintext[12]), .B(
        Red_RoundKey[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_1_U1 ( .A(Red_Plaintext[13]), .B(
        Red_RoundKey[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_2_U1 ( .A(Red_Plaintext[14]), .B(
        Red_RoundKey[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_0_U1 ( .A(Red_Plaintext[15]), .B(
        Red_RoundKey[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_1_U1 ( .A(Red_Plaintext[16]), .B(
        Red_RoundKey[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_2_U1 ( .A(Red_Plaintext[17]), .B(
        Red_RoundKey[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_0_U1 ( .A(Red_Plaintext[18]), .B(
        Red_RoundKey[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_1_U1 ( .A(Red_Plaintext[19]), .B(
        Red_RoundKey[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_2_U1 ( .A(Red_Plaintext[20]), .B(
        Red_RoundKey[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_0_U1 ( .A(Red_Plaintext[21]), .B(
        Red_RoundKey[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_1_U1 ( .A(Red_Plaintext[22]), .B(
        Red_RoundKey[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_2_U1 ( .A(Red_Plaintext[23]), .B(
        Red_RoundKey[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_0_U1 ( .A(Red_Plaintext[24]), .B(
        Red_RoundKey[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_1_U1 ( .A(Red_Plaintext[25]), .B(
        Red_RoundKey[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_2_U1 ( .A(Red_Plaintext[26]), .B(
        Red_RoundKey[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_0_U1 ( .A(Red_Plaintext[27]), .B(
        Red_RoundKey[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_1_U1 ( .A(Red_Plaintext[28]), .B(
        Red_RoundKey[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_2_U1 ( .A(Red_Plaintext[29]), .B(
        Red_RoundKey[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_0_U1 ( .A(Red_Plaintext[30]), .B(
        Red_RoundKey[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_1_U1 ( .A(Red_Plaintext[31]), .B(
        Red_RoundKey[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_2_U1 ( .A(Red_Plaintext[32]), .B(
        Red_RoundKey[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_0_U1 ( .A(Red_Plaintext[33]), .B(
        Red_RoundKey[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_1_U1 ( .A(Red_Plaintext[34]), .B(
        Red_RoundKey[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_2_U1 ( .A(Red_Plaintext[35]), .B(
        Red_RoundKey[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_0_U1 ( .A(Red_Plaintext[36]), .B(
        Red_RoundKey[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_1_U1 ( .A(Red_Plaintext[37]), .B(
        Red_RoundKey[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_2_U1 ( .A(Red_Plaintext[38]), .B(
        Red_RoundKey[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_0_U1 ( .A(Red_Plaintext[39]), .B(
        Red_RoundKey[39]), .Z(Red_AddRoundKeyOutput[39]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_1_U1 ( .A(Red_Plaintext[40]), .B(
        Red_RoundKey[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_2_U1 ( .A(Red_Plaintext[41]), .B(
        Red_RoundKey[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_0_U1 ( .A(Red_Plaintext[42]), .B(
        Red_RoundKey[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_1_U1 ( .A(Red_Plaintext[43]), .B(
        Red_RoundKey[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_2_U1 ( .A(Red_Plaintext[44]), .B(
        Red_RoundKey[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_0_U1 ( .A(Red_Plaintext[45]), .B(
        Red_RoundKey[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_1_U1 ( .A(Red_Plaintext[46]), .B(
        Red_RoundKey[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_2_U1 ( .A(Red_Plaintext[47]), .B(
        Red_RoundKey[47]), .Z(Red_AddRoundKeyOutput[47]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[9]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U4 ( .A1(AddRoundKeyOutput[2]), 
        .A2(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U3 ( .A1(AddRoundKeyOutput[0]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U2 ( .A1(AddRoundKeyOutput[2]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput[1]), 
        .B(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_0_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[10]) );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U2 ( .A1(AddRoundKeyOutput[3]), 
        .A2(AddRoundKeyOutput[2]), .ZN(Red_SubCellInst_LFInst_0_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U1 ( .A1(AddRoundKeyOutput[1]), 
        .A2(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_0_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[11])
         );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(AddRoundKeyOutput[1]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U4 ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[0]), .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n13), .A2(AddRoundKeyOutput[3]), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n12), .A2(AddRoundKeyOutput[2]), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U1 ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[0]) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U4 ( .A1(AddRoundKeyOutput[6]), 
        .A2(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U3 ( .A1(AddRoundKeyOutput[4]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U2 ( .A1(AddRoundKeyOutput[6]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput[5]), 
        .B(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_1_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[1]) );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U2 ( .A1(AddRoundKeyOutput[7]), 
        .A2(AddRoundKeyOutput[6]), .ZN(Red_SubCellInst_LFInst_1_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U1 ( .A1(AddRoundKeyOutput[5]), 
        .A2(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n16), .A2(
        Red_SubCellInst_LFInst_1_LFInst_2_n15), .ZN(Red_ShiftRowsOutput[2]) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n14), .A2(AddRoundKeyOutput[7]), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U4 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n13), .A2(AddRoundKeyOutput[6]), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U3 ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n13)
         );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U2 ( .A1(AddRoundKeyOutput[5]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[4]), .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[3]) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U4 ( .A1(AddRoundKeyOutput[10]), 
        .A2(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U3 ( .A1(AddRoundKeyOutput[8]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U2 ( .A1(AddRoundKeyOutput[10]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput[9]), 
        .B(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_2_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[4]) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U2 ( .A1(AddRoundKeyOutput[11]), 
        .A2(AddRoundKeyOutput[10]), .ZN(Red_SubCellInst_LFInst_2_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U1 ( .A1(AddRoundKeyOutput[9]), 
        .A2(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_2_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[5]) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(AddRoundKeyOutput[9]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U4 ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[8]), .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n13), .A2(AddRoundKeyOutput[11]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n12), .A2(AddRoundKeyOutput[10]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U1 ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[6]) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U4 ( .A1(AddRoundKeyOutput[14]), 
        .A2(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U3 ( .A1(AddRoundKeyOutput[12]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U2 ( .A1(AddRoundKeyOutput[14]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput[13]), 
        .B(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_3_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[7]) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U2 ( .A1(AddRoundKeyOutput[15]), 
        .A2(AddRoundKeyOutput[14]), .ZN(Red_SubCellInst_LFInst_3_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U1 ( .A1(AddRoundKeyOutput[13]), 
        .A2(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_3_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[8]) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(AddRoundKeyOutput[13]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U4 ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[12]), .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n13), .A2(AddRoundKeyOutput[15]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n12), .A2(AddRoundKeyOutput[14]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U1 ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_4_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[18])
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U4 ( .A1(AddRoundKeyOutput[18]), 
        .A2(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(AddRoundKeyOutput[16]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U2 ( .A1(AddRoundKeyOutput[18]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[17]), 
        .B(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_4_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[19]) );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U2 ( .A1(AddRoundKeyOutput[19]), 
        .A2(AddRoundKeyOutput[18]), .ZN(Red_SubCellInst_LFInst_4_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(AddRoundKeyOutput[17]), 
        .A2(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_4_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[20])
         );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U5 ( .A1(AddRoundKeyOutput[17]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U4 ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[16]), .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n13), .A2(AddRoundKeyOutput[19]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n12), .A2(AddRoundKeyOutput[18]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U1 ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_5_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[21])
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U4 ( .A1(AddRoundKeyOutput[22]), 
        .A2(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(AddRoundKeyOutput[20]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U2 ( .A1(AddRoundKeyOutput[22]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[21]), 
        .B(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_5_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[22]) );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U2 ( .A1(AddRoundKeyOutput[23]), 
        .A2(AddRoundKeyOutput[22]), .ZN(Red_SubCellInst_LFInst_5_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(AddRoundKeyOutput[21]), 
        .A2(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_5_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[23])
         );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U5 ( .A1(AddRoundKeyOutput[21]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U4 ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[20]), .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n13), .A2(AddRoundKeyOutput[23]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n12), .A2(AddRoundKeyOutput[22]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U1 ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_6_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[12])
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U4 ( .A1(AddRoundKeyOutput[26]), 
        .A2(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(AddRoundKeyOutput[24]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U2 ( .A1(AddRoundKeyOutput[26]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[25]), 
        .B(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_6_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[13]) );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U2 ( .A1(AddRoundKeyOutput[27]), 
        .A2(AddRoundKeyOutput[26]), .ZN(Red_SubCellInst_LFInst_6_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(AddRoundKeyOutput[25]), 
        .A2(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U7 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n17), .A2(
        Red_SubCellInst_LFInst_6_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[14])
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n15), .A2(AddRoundKeyOutput[27]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n14), .A2(AddRoundKeyOutput[26]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U4 ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n13), .A2(
        Red_SubCellInst_LFInst_6_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_2_n17) );
  INV_X1 Red_SubCellInst_LFInst_6_LFInst_2_U2 ( .A(AddRoundKeyOutput[25]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[26]), .Z(Red_SubCellInst_LFInst_6_LFInst_2_n13)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_7_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[15])
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U4 ( .A1(AddRoundKeyOutput[30]), 
        .A2(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(AddRoundKeyOutput[28]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U2 ( .A1(AddRoundKeyOutput[30]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[29]), 
        .B(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_7_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[16]) );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U2 ( .A1(AddRoundKeyOutput[31]), 
        .A2(AddRoundKeyOutput[30]), .ZN(Red_SubCellInst_LFInst_7_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(AddRoundKeyOutput[29]), 
        .A2(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_7_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[17])
         );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U5 ( .A1(AddRoundKeyOutput[29]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U4 ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[28]), .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n13), .A2(AddRoundKeyOutput[31]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n12), .A2(AddRoundKeyOutput[30]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U1 ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[27])
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U4 ( .A1(AddRoundKeyOutput[34]), 
        .A2(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U3 ( .A1(AddRoundKeyOutput[32]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U2 ( .A1(AddRoundKeyOutput[34]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput[33]), 
        .B(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_8_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[28]) );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(AddRoundKeyOutput[35]), 
        .A2(AddRoundKeyOutput[34]), .ZN(Red_SubCellInst_LFInst_8_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U1 ( .A1(AddRoundKeyOutput[33]), 
        .A2(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n11), .A2(
        Red_SubCellInst_LFInst_8_LFInst_2_n13), .ZN(Red_ShiftRowsOutput[29])
         );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U5 ( .A1(AddRoundKeyOutput[33]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_2_n13) );
  XNOR2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U4 ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[32]), .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n10), .A2(AddRoundKeyOutput[35]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n11) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n9), .A2(AddRoundKeyOutput[34]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n10) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U1 ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[30])
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U4 ( .A1(AddRoundKeyOutput[38]), 
        .A2(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U3 ( .A1(AddRoundKeyOutput[36]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U2 ( .A1(AddRoundKeyOutput[38]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput[37]), 
        .B(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_9_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[31]) );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(AddRoundKeyOutput[39]), 
        .A2(AddRoundKeyOutput[38]), .ZN(Red_SubCellInst_LFInst_9_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U1 ( .A1(AddRoundKeyOutput[37]), 
        .A2(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_9_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[32])
         );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(AddRoundKeyOutput[37]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U4 ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[36]), .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n13), .A2(AddRoundKeyOutput[39]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n12), .A2(AddRoundKeyOutput[38]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U1 ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[33])
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U4 ( .A1(AddRoundKeyOutput[42]), 
        .A2(AddRoundKeyOutput[43]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U3 ( .A1(AddRoundKeyOutput[40]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U2 ( .A1(AddRoundKeyOutput[42]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput[41]), 
        .B(AddRoundKeyOutput[43]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_10_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[34])
         );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(AddRoundKeyOutput[43]), 
        .A2(AddRoundKeyOutput[42]), .ZN(Red_SubCellInst_LFInst_10_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U1 ( .A1(AddRoundKeyOutput[41]), 
        .A2(AddRoundKeyOutput[43]), .ZN(Red_SubCellInst_LFInst_10_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_10_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[35])
         );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(AddRoundKeyOutput[41]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U4 ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[40]), .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n13), .A2(AddRoundKeyOutput[43]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n12), .A2(AddRoundKeyOutput[42]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U1 ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[24])
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U4 ( .A1(AddRoundKeyOutput[46]), 
        .A2(AddRoundKeyOutput[47]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U3 ( .A1(AddRoundKeyOutput[44]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U2 ( .A1(AddRoundKeyOutput[46]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput[45]), 
        .B(AddRoundKeyOutput[47]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_11_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[25])
         );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(AddRoundKeyOutput[47]), 
        .A2(AddRoundKeyOutput[46]), .ZN(Red_SubCellInst_LFInst_11_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U1 ( .A1(AddRoundKeyOutput[45]), 
        .A2(AddRoundKeyOutput[47]), .ZN(Red_SubCellInst_LFInst_11_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_11_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[26])
         );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(AddRoundKeyOutput[45]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U4 ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[44]), .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n13), .A2(AddRoundKeyOutput[47]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n12), .A2(AddRoundKeyOutput[46]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U1 ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[36])
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U4 ( .A1(AddRoundKeyOutput[50]), 
        .A2(AddRoundKeyOutput[51]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U3 ( .A1(AddRoundKeyOutput[48]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U2 ( .A1(AddRoundKeyOutput[50]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput[49]), 
        .B(AddRoundKeyOutput[51]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_12_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[37])
         );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U2 ( .A1(AddRoundKeyOutput[51]), 
        .A2(AddRoundKeyOutput[50]), .ZN(Red_SubCellInst_LFInst_12_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U1 ( .A1(AddRoundKeyOutput[49]), 
        .A2(AddRoundKeyOutput[51]), .ZN(Red_SubCellInst_LFInst_12_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_12_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[38])
         );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U5 ( .A1(AddRoundKeyOutput[49]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U4 ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[48]), .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n13), .A2(AddRoundKeyOutput[51]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n12), .A2(AddRoundKeyOutput[50]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U1 ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[39])
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U4 ( .A1(AddRoundKeyOutput[54]), 
        .A2(AddRoundKeyOutput[55]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U2 ( .A1(AddRoundKeyOutput[54]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput[53]), 
        .B(AddRoundKeyOutput[55]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_13_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[40])
         );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U2 ( .A1(AddRoundKeyOutput[55]), 
        .A2(AddRoundKeyOutput[54]), .ZN(Red_SubCellInst_LFInst_13_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U1 ( .A1(AddRoundKeyOutput[53]), 
        .A2(AddRoundKeyOutput[55]), .ZN(Red_SubCellInst_LFInst_13_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n16), .A2(
        Red_SubCellInst_LFInst_13_LFInst_2_n15), .ZN(Red_ShiftRowsOutput[41])
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U5 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n14), .A2(AddRoundKeyOutput[55]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U4 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n13), .A2(AddRoundKeyOutput[54]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U3 ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n13) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U2 ( .A1(AddRoundKeyOutput[53]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_2_n12), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[52]), .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n12)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[42])
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U4 ( .A1(AddRoundKeyOutput[58]), 
        .A2(AddRoundKeyOutput[59]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U3 ( .A1(AddRoundKeyOutput[56]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U2 ( .A1(AddRoundKeyOutput[58]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput[57]), 
        .B(AddRoundKeyOutput[59]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_14_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[43])
         );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U2 ( .A1(AddRoundKeyOutput[59]), 
        .A2(AddRoundKeyOutput[58]), .ZN(Red_SubCellInst_LFInst_14_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U1 ( .A1(AddRoundKeyOutput[57]), 
        .A2(AddRoundKeyOutput[59]), .ZN(Red_SubCellInst_LFInst_14_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_14_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[44])
         );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U5 ( .A1(AddRoundKeyOutput[57]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U4 ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[56]), .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n13), .A2(AddRoundKeyOutput[59]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n12), .A2(AddRoundKeyOutput[58]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U1 ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n12), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n11), .ZN(Red_ShiftRowsOutput[45])
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U4 ( .A1(AddRoundKeyOutput[62]), 
        .A2(AddRoundKeyOutput[63]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U3 ( .A1(AddRoundKeyOutput[60]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_0_n10), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U2 ( .A1(AddRoundKeyOutput[62]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_0_n9), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput[61]), 
        .B(AddRoundKeyOutput[63]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n9)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U3 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_1_n6), .A2(
        Red_SubCellInst_LFInst_15_LFInst_1_n5), .ZN(Red_ShiftRowsOutput[46])
         );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U2 ( .A1(AddRoundKeyOutput[63]), 
        .A2(AddRoundKeyOutput[62]), .ZN(Red_SubCellInst_LFInst_15_LFInst_1_n5)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U1 ( .A1(AddRoundKeyOutput[61]), 
        .A2(AddRoundKeyOutput[63]), .ZN(Red_SubCellInst_LFInst_15_LFInst_1_n6)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n14), .A2(
        Red_SubCellInst_LFInst_15_LFInst_2_n16), .ZN(Red_ShiftRowsOutput[47])
         );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U5 ( .A1(AddRoundKeyOutput[61]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_2_n15), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U4 ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[60]), .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n15)
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U3 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n13), .A2(AddRoundKeyOutput[63]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U2 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n12), .A2(AddRoundKeyOutput[62]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U1 ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n12) );
  BUF_X1 Red_MCInst_MC0_U3 ( .A(ShiftRowsOutput[28]), .Z(
        Red_MCInst_MC0_v2_1[1]) );
  BUF_X1 Red_MCInst_MC0_U2 ( .A(MCInst_MC0_v1_3[2]), .Z(Red_MCInst_MC0_v1_2[1]) );
  XOR2_X1 Red_MCInst_MC0_v0_2Inst_0_U1 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(Red_MCInst_MC0_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC0_v0_3Inst_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U2 ( .A(Red_MCInst_MC0_v1_0Inst_0_n3), 
        .B(MCInst_MC0_v1_3[3]), .ZN(Red_MCInst_MC0_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC0_v1_2Inst_0_U1 ( .A(Red_MCInst_MC0_v1_2[1]), .B(
        Red_MCInst_MC0_v1_1[2]), .Z(Red_MCInst_MC0_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC0_v1_3Inst_0_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .Z(Red_MCInst_MC0_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC0_v2_0Inst_0_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(Red_MCInst_MC0_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC0_v2_1Inst_0_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC0_v2_2Inst_0_U2 ( .A(Red_MCInst_MC0_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC0_v2_2[1]), .ZN(Red_MCInst_MC0_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC0_v2_2Inst_0_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[2]), .ZN(Red_MCInst_MC0_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC0_v2_3Inst_0_U2 ( .A(Red_MCInst_MC0_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC0_v2_2[1]), .ZN(Red_MCInst_MC0_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC0_v2_3Inst_0_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[3]), .ZN(Red_MCInst_MC0_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC0_v3_0Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U3 ( .A(Red_MCInst_MC0_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC0_v3_2Inst_0_n5), .ZN(Red_MCInst_MC0_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U2 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC0_v3_3Inst_0_U1 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .Z(Red_MCInst_MC0_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC0_v0_0Inst_1_U1 ( .A(Red_MCInst_MC0_v0_2[2]), .B(
        Red_MCInst_MC0_v0_1[0]), .Z(Red_MCInst_MC0_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC0_v0_1Inst_1_U2 ( .A(Red_MCInst_MC0_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC0_v0_1[0]), .ZN(Red_MCInst_MC0_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC0_v0_1Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .ZN(Red_MCInst_MC0_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        MCInst_MC0_v0_3[3]), .Z(Red_MCInst_MC0_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_1_U2 ( .A(Red_MCInst_MC0_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_1Inst_1_U3 ( .A(Red_MCInst_MC0_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC0_v1_1Inst_1_n5), .ZN(Red_MCInst_MC0_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC0_v1_1Inst_1_U2 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC0_v1_1Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .Z(Red_MCInst_MC0_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC0_v1_3Inst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[3]), .Z(Red_MCInst_MC0_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC0_v2_0Inst_1_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC0_v2_3Inst_1_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(Red_MCInst_MC0_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC0_v3_0Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .Z(Red_MCInst_MC0_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC0_v3_1Inst_1_U3 ( .A(Red_MCInst_MC0_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC0_v3_1Inst_1_n5), .ZN(Red_MCInst_MC0_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC0_v3_1Inst_1_U2 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC0_v3_1Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC0_v3_2Inst_1_U1 ( .A(Red_MCInst_MC0_v3_3[2]), .B(
        MCInst_MC0_v3_0[3]), .Z(Red_MCInst_MC0_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC0_v3_3Inst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC0_v0_0Inst_2_U2 ( .A(Red_MCInst_MC0_v0_0Inst_2_n3), 
        .B(MCInst_MC0_v0_3[3]), .ZN(Red_MCInst_MC0_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .ZN(Red_MCInst_MC0_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC0_v0_1Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_2_U3 ( .A(Red_MCInst_MC0_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC0_v0_3Inst_2_n5), .ZN(Red_MCInst_MC0_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_2_U2 ( .A(MCInst_MC0_v0_3[3]), .B(
        Red_MCInst_MC0_v0_1[0]), .ZN(Red_MCInst_MC0_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v0_3Inst_2_U1 ( .A(Red_MCInst_MC0_v0_0[0]), .B(
        Red_MCInst_MC0_v0_2[2]), .Z(Red_MCInst_MC0_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_2_U2 ( .A(Red_MCInst_MC0_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_2_U1 ( .A(Red_MCInst_MC0_v1_2[1]), .B(
        MCInst_MC0_v1_3[3]), .ZN(Red_MCInst_MC0_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_2Inst_2_U2 ( .A(Red_MCInst_MC0_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC0_v1_2Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_2_U3 ( .A(Red_MCInst_MC0_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC0_v1_3Inst_2_n5), .ZN(Red_MCInst_MC0_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_2_U2 ( .A(MCInst_MC0_v1_3[3]), .B(
        Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v1_3Inst_2_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        Red_MCInst_MC0_v1_2[1]), .Z(Red_MCInst_MC0_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_2_U3 ( .A(Red_MCInst_MC0_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC0_v2_0Inst_2_n5), .ZN(Red_MCInst_MC0_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_2_U2 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .ZN(Red_MCInst_MC0_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v2_0Inst_2_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[2]), .Z(Red_MCInst_MC0_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC0_v2_1Inst_2_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(Red_MCInst_MC0_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC0_v2_2Inst_2_U1 ( .A(MCInst_MC0_v2_0[3]), .B(
        Red_MCInst_MC0_v2_2[1]), .Z(Red_MCInst_MC0_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC0_v2_3Inst_2_U1 ( .A(Red_MCInst_MC0_v2_1[1]), .B(
        MCInst_MC0_v2_0[3]), .Z(Red_MCInst_MC0_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_2_U3 ( .A(Red_MCInst_MC0_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC0_v3_0Inst_2_n5), .ZN(Red_MCInst_MC0_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_2_U2 ( .A(MCInst_MC0_v3_0[3]), .B(
        Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC0_v3_0Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_2_U2 ( .A(Red_MCInst_MC0_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC0_v3_1[2]), .ZN(Red_MCInst_MC0_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_2_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        MCInst_MC0_v3_0[3]), .ZN(Red_MCInst_MC0_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[45]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_0[0]), 
        .B(Red_MCInst_MC0_v1_0[0]), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), 
        .B(Red_MCInst_MC0_v3_0[0]), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[46]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_0[1]), 
        .B(Red_MCInst_MC0_v1_0[1]), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_0[1]), 
        .B(Red_MCInst_MC0_v3_0[1]), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[47]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_0[2]), 
        .B(Red_MCInst_MC0_v1_0[2]), .ZN(Red_MCInst_MC0_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_0[2]), 
        .B(Red_MCInst_MC0_v3_0[2]), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[33]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_1[0]), 
        .B(Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_1[0]), 
        .B(Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[34]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_1[1]), 
        .B(Red_MCInst_MC0_v1_1[1]), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_1[1]), 
        .B(Red_MCInst_MC0_v3_1[1]), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[35]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_1[2]), 
        .B(Red_MCInst_MC0_v1_1[2]), .ZN(Red_MCInst_MC0_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_1[2]), 
        .B(Red_MCInst_MC0_v3_1[2]), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[21]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_2[0]), 
        .B(Red_MCInst_MC0_v1_2[0]), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_2[0]), 
        .B(Red_MCInst_MC0_v3_2[0]), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[22]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_2[1]), 
        .B(Red_MCInst_MC0_v1_2[1]), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_2[1]), 
        .B(Red_MCInst_MC0_v3_2[1]), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[23]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_2[2]), 
        .B(Red_MCInst_MC0_v1_2[2]), .ZN(Red_MCInst_MC0_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), 
        .B(Red_MCInst_MC0_v3_2[2]), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[9]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC0_v2_3[0]), 
        .B(Red_MCInst_MC0_v1_3[0]), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC0_v0_3[0]), 
        .B(Red_MCInst_MC0_v3_3[0]), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[10]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC0_v2_3[1]), 
        .B(Red_MCInst_MC0_v1_3[1]), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC0_v0_3[1]), 
        .B(Red_MCInst_MC0_v3_3[1]), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[11]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC0_v2_3[2]), 
        .B(Red_MCInst_MC0_v1_3[2]), .ZN(Red_MCInst_MC0_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC0_v0_3[2]), 
        .B(Red_MCInst_MC0_v3_3[2]), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst_MC1_U3 ( .A(ShiftRowsOutput[24]), .Z(
        Red_MCInst_MC1_v2_1[1]) );
  BUF_X1 Red_MCInst_MC1_U2 ( .A(MCInst_MC1_v1_3[2]), .Z(Red_MCInst_MC1_v1_2[1]) );
  XOR2_X1 Red_MCInst_MC1_v0_2Inst_0_U1 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(Red_MCInst_MC1_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC1_v0_3Inst_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U2 ( .A(Red_MCInst_MC1_v1_0Inst_0_n3), 
        .B(MCInst_MC1_v1_3[3]), .ZN(Red_MCInst_MC1_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC1_v1_2Inst_0_U1 ( .A(Red_MCInst_MC1_v1_2[1]), .B(
        Red_MCInst_MC1_v1_1[2]), .Z(Red_MCInst_MC1_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC1_v1_3Inst_0_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .Z(Red_MCInst_MC1_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC1_v2_0Inst_0_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(Red_MCInst_MC1_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC1_v2_1Inst_0_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC1_v2_2Inst_0_U2 ( .A(Red_MCInst_MC1_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC1_v2_2[1]), .ZN(Red_MCInst_MC1_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC1_v2_2Inst_0_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[2]), .ZN(Red_MCInst_MC1_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC1_v2_3Inst_0_U2 ( .A(Red_MCInst_MC1_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC1_v2_2[1]), .ZN(Red_MCInst_MC1_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC1_v2_3Inst_0_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[3]), .ZN(Red_MCInst_MC1_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC1_v3_0Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U3 ( .A(Red_MCInst_MC1_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC1_v3_2Inst_0_n5), .ZN(Red_MCInst_MC1_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U2 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC1_v3_3Inst_0_U1 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .Z(Red_MCInst_MC1_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC1_v0_0Inst_1_U1 ( .A(Red_MCInst_MC1_v0_2[2]), .B(
        Red_MCInst_MC1_v0_1[0]), .Z(Red_MCInst_MC1_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC1_v0_1Inst_1_U2 ( .A(Red_MCInst_MC1_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC1_v0_1[0]), .ZN(Red_MCInst_MC1_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC1_v0_1Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .ZN(Red_MCInst_MC1_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        MCInst_MC1_v0_3[3]), .Z(Red_MCInst_MC1_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_1_U2 ( .A(Red_MCInst_MC1_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_1Inst_1_U3 ( .A(Red_MCInst_MC1_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC1_v1_1Inst_1_n5), .ZN(Red_MCInst_MC1_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC1_v1_1Inst_1_U2 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC1_v1_1Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .Z(Red_MCInst_MC1_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC1_v1_3Inst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[3]), .Z(Red_MCInst_MC1_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC1_v2_0Inst_1_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC1_v2_3Inst_1_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(Red_MCInst_MC1_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC1_v3_0Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .Z(Red_MCInst_MC1_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC1_v3_1Inst_1_U3 ( .A(Red_MCInst_MC1_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC1_v3_1Inst_1_n5), .ZN(Red_MCInst_MC1_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC1_v3_1Inst_1_U2 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC1_v3_1Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC1_v3_2Inst_1_U1 ( .A(Red_MCInst_MC1_v3_3[2]), .B(
        MCInst_MC1_v3_0[3]), .Z(Red_MCInst_MC1_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC1_v3_3Inst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC1_v0_0Inst_2_U2 ( .A(Red_MCInst_MC1_v0_0Inst_2_n3), 
        .B(MCInst_MC1_v0_3[3]), .ZN(Red_MCInst_MC1_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .ZN(Red_MCInst_MC1_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC1_v0_1Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_2_U3 ( .A(Red_MCInst_MC1_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC1_v0_3Inst_2_n5), .ZN(Red_MCInst_MC1_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_2_U2 ( .A(MCInst_MC1_v0_3[3]), .B(
        Red_MCInst_MC1_v0_1[0]), .ZN(Red_MCInst_MC1_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v0_3Inst_2_U1 ( .A(Red_MCInst_MC1_v0_0[0]), .B(
        Red_MCInst_MC1_v0_2[2]), .Z(Red_MCInst_MC1_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_2_U2 ( .A(Red_MCInst_MC1_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_2_U1 ( .A(Red_MCInst_MC1_v1_2[1]), .B(
        MCInst_MC1_v1_3[3]), .ZN(Red_MCInst_MC1_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_2Inst_2_U2 ( .A(Red_MCInst_MC1_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC1_v1_2Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_2_U3 ( .A(Red_MCInst_MC1_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC1_v1_3Inst_2_n5), .ZN(Red_MCInst_MC1_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_2_U2 ( .A(MCInst_MC1_v1_3[3]), .B(
        Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v1_3Inst_2_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        Red_MCInst_MC1_v1_2[1]), .Z(Red_MCInst_MC1_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_2_U3 ( .A(Red_MCInst_MC1_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC1_v2_0Inst_2_n5), .ZN(Red_MCInst_MC1_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_2_U2 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .ZN(Red_MCInst_MC1_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v2_0Inst_2_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[2]), .Z(Red_MCInst_MC1_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC1_v2_1Inst_2_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(Red_MCInst_MC1_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC1_v2_2Inst_2_U1 ( .A(MCInst_MC1_v2_0[3]), .B(
        Red_MCInst_MC1_v2_2[1]), .Z(Red_MCInst_MC1_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC1_v2_3Inst_2_U1 ( .A(Red_MCInst_MC1_v2_1[1]), .B(
        MCInst_MC1_v2_0[3]), .Z(Red_MCInst_MC1_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_2_U3 ( .A(Red_MCInst_MC1_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC1_v3_0Inst_2_n5), .ZN(Red_MCInst_MC1_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_2_U2 ( .A(MCInst_MC1_v3_0[3]), .B(
        Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC1_v3_0Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_2_U2 ( .A(Red_MCInst_MC1_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC1_v3_1[2]), .ZN(Red_MCInst_MC1_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_2_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        MCInst_MC1_v3_0[3]), .ZN(Red_MCInst_MC1_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[42]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_0[0]), 
        .B(Red_MCInst_MC1_v1_0[0]), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), 
        .B(Red_MCInst_MC1_v3_0[0]), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[43]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_0[1]), 
        .B(Red_MCInst_MC1_v1_0[1]), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_0[1]), 
        .B(Red_MCInst_MC1_v3_0[1]), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[44]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_0[2]), 
        .B(Red_MCInst_MC1_v1_0[2]), .ZN(Red_MCInst_MC1_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_0[2]), 
        .B(Red_MCInst_MC1_v3_0[2]), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[30]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_1[0]), 
        .B(Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_1[0]), 
        .B(Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[31]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_1[1]), 
        .B(Red_MCInst_MC1_v1_1[1]), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_1[1]), 
        .B(Red_MCInst_MC1_v3_1[1]), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[32]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_1[2]), 
        .B(Red_MCInst_MC1_v1_1[2]), .ZN(Red_MCInst_MC1_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_1[2]), 
        .B(Red_MCInst_MC1_v3_1[2]), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[18]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_2[0]), 
        .B(Red_MCInst_MC1_v1_2[0]), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_2[0]), 
        .B(Red_MCInst_MC1_v3_2[0]), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[19]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_2[1]), 
        .B(Red_MCInst_MC1_v1_2[1]), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_2[1]), 
        .B(Red_MCInst_MC1_v3_2[1]), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[20]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_2[2]), 
        .B(Red_MCInst_MC1_v1_2[2]), .ZN(Red_MCInst_MC1_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), 
        .B(Red_MCInst_MC1_v3_2[2]), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[6]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC1_v2_3[0]), 
        .B(Red_MCInst_MC1_v1_3[0]), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC1_v0_3[0]), 
        .B(Red_MCInst_MC1_v3_3[0]), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[7]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC1_v2_3[1]), 
        .B(Red_MCInst_MC1_v1_3[1]), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC1_v0_3[1]), 
        .B(Red_MCInst_MC1_v3_3[1]), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[8]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC1_v2_3[2]), 
        .B(Red_MCInst_MC1_v1_3[2]), .ZN(Red_MCInst_MC1_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC1_v0_3[2]), 
        .B(Red_MCInst_MC1_v3_3[2]), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst_MC2_U3 ( .A(ShiftRowsOutput[20]), .Z(
        Red_MCInst_MC2_v2_1[1]) );
  BUF_X1 Red_MCInst_MC2_U2 ( .A(MCInst_MC2_v1_3[2]), .Z(Red_MCInst_MC2_v1_2[1]) );
  XOR2_X1 Red_MCInst_MC2_v0_2Inst_0_U1 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(Red_MCInst_MC2_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC2_v0_3Inst_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U2 ( .A(Red_MCInst_MC2_v1_0Inst_0_n3), 
        .B(MCInst_MC2_v1_3[3]), .ZN(Red_MCInst_MC2_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC2_v1_2Inst_0_U1 ( .A(Red_MCInst_MC2_v1_2[1]), .B(
        Red_MCInst_MC2_v1_1[2]), .Z(Red_MCInst_MC2_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC2_v1_3Inst_0_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .Z(Red_MCInst_MC2_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC2_v2_0Inst_0_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(Red_MCInst_MC2_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC2_v2_1Inst_0_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC2_v2_2Inst_0_U2 ( .A(Red_MCInst_MC2_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC2_v2_2[1]), .ZN(Red_MCInst_MC2_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC2_v2_2Inst_0_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[2]), .ZN(Red_MCInst_MC2_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC2_v2_3Inst_0_U2 ( .A(Red_MCInst_MC2_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC2_v2_2[1]), .ZN(Red_MCInst_MC2_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC2_v2_3Inst_0_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[3]), .ZN(Red_MCInst_MC2_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC2_v3_0Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U3 ( .A(Red_MCInst_MC2_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC2_v3_2Inst_0_n5), .ZN(Red_MCInst_MC2_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U2 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC2_v3_3Inst_0_U1 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .Z(Red_MCInst_MC2_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC2_v0_0Inst_1_U1 ( .A(Red_MCInst_MC2_v0_2[2]), .B(
        Red_MCInst_MC2_v0_1[0]), .Z(Red_MCInst_MC2_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC2_v0_1Inst_1_U2 ( .A(Red_MCInst_MC2_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC2_v0_1[0]), .ZN(Red_MCInst_MC2_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC2_v0_1Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .ZN(Red_MCInst_MC2_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        MCInst_MC2_v0_3[3]), .Z(Red_MCInst_MC2_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_1_U2 ( .A(Red_MCInst_MC2_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_1Inst_1_U3 ( .A(Red_MCInst_MC2_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC2_v1_1Inst_1_n5), .ZN(Red_MCInst_MC2_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC2_v1_1Inst_1_U2 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC2_v1_1Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .Z(Red_MCInst_MC2_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC2_v1_3Inst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[3]), .Z(Red_MCInst_MC2_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC2_v2_0Inst_1_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC2_v2_3Inst_1_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(Red_MCInst_MC2_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC2_v3_0Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .Z(Red_MCInst_MC2_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC2_v3_1Inst_1_U3 ( .A(Red_MCInst_MC2_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC2_v3_1Inst_1_n5), .ZN(Red_MCInst_MC2_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC2_v3_1Inst_1_U2 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC2_v3_1Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC2_v3_2Inst_1_U1 ( .A(Red_MCInst_MC2_v3_3[2]), .B(
        MCInst_MC2_v3_0[3]), .Z(Red_MCInst_MC2_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC2_v3_3Inst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC2_v0_0Inst_2_U2 ( .A(Red_MCInst_MC2_v0_0Inst_2_n3), 
        .B(MCInst_MC2_v0_3[3]), .ZN(Red_MCInst_MC2_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .ZN(Red_MCInst_MC2_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC2_v0_1Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_2_U3 ( .A(Red_MCInst_MC2_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC2_v0_3Inst_2_n5), .ZN(Red_MCInst_MC2_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_2_U2 ( .A(MCInst_MC2_v0_3[3]), .B(
        Red_MCInst_MC2_v0_1[0]), .ZN(Red_MCInst_MC2_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v0_3Inst_2_U1 ( .A(Red_MCInst_MC2_v0_0[0]), .B(
        Red_MCInst_MC2_v0_2[2]), .Z(Red_MCInst_MC2_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_2_U2 ( .A(Red_MCInst_MC2_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_2_U1 ( .A(Red_MCInst_MC2_v1_2[1]), .B(
        MCInst_MC2_v1_3[3]), .ZN(Red_MCInst_MC2_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_2Inst_2_U2 ( .A(Red_MCInst_MC2_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC2_v1_2Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_2_U3 ( .A(Red_MCInst_MC2_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC2_v1_3Inst_2_n5), .ZN(Red_MCInst_MC2_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_2_U2 ( .A(MCInst_MC2_v1_3[3]), .B(
        Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v1_3Inst_2_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        Red_MCInst_MC2_v1_2[1]), .Z(Red_MCInst_MC2_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_2_U3 ( .A(Red_MCInst_MC2_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC2_v2_0Inst_2_n5), .ZN(Red_MCInst_MC2_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_2_U2 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .ZN(Red_MCInst_MC2_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v2_0Inst_2_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[2]), .Z(Red_MCInst_MC2_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC2_v2_1Inst_2_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(Red_MCInst_MC2_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC2_v2_2Inst_2_U1 ( .A(MCInst_MC2_v2_0[3]), .B(
        Red_MCInst_MC2_v2_2[1]), .Z(Red_MCInst_MC2_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC2_v2_3Inst_2_U1 ( .A(Red_MCInst_MC2_v2_1[1]), .B(
        MCInst_MC2_v2_0[3]), .Z(Red_MCInst_MC2_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_2_U3 ( .A(Red_MCInst_MC2_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC2_v3_0Inst_2_n5), .ZN(Red_MCInst_MC2_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_2_U2 ( .A(MCInst_MC2_v3_0[3]), .B(
        Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC2_v3_0Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_2_U2 ( .A(Red_MCInst_MC2_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC2_v3_1[2]), .ZN(Red_MCInst_MC2_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_2_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        MCInst_MC2_v3_0[3]), .ZN(Red_MCInst_MC2_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[39]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_0[0]), 
        .B(Red_MCInst_MC2_v1_0[0]), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), 
        .B(Red_MCInst_MC2_v3_0[0]), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[40]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_0[1]), 
        .B(Red_MCInst_MC2_v1_0[1]), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_0[1]), 
        .B(Red_MCInst_MC2_v3_0[1]), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[41]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_0[2]), 
        .B(Red_MCInst_MC2_v1_0[2]), .ZN(Red_MCInst_MC2_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_0[2]), 
        .B(Red_MCInst_MC2_v3_0[2]), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[27]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_1[0]), 
        .B(Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_1[0]), 
        .B(Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[28]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_1[1]), 
        .B(Red_MCInst_MC2_v1_1[1]), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_1[1]), 
        .B(Red_MCInst_MC2_v3_1[1]), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[29]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_1[2]), 
        .B(Red_MCInst_MC2_v1_1[2]), .ZN(Red_MCInst_MC2_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_1[2]), 
        .B(Red_MCInst_MC2_v3_1[2]), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[15]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_2[0]), 
        .B(Red_MCInst_MC2_v1_2[0]), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_2[0]), 
        .B(Red_MCInst_MC2_v3_2[0]), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[16]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_2[1]), 
        .B(Red_MCInst_MC2_v1_2[1]), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_2[1]), 
        .B(Red_MCInst_MC2_v3_2[1]), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[17]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_2[2]), 
        .B(Red_MCInst_MC2_v1_2[2]), .ZN(Red_MCInst_MC2_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), 
        .B(Red_MCInst_MC2_v3_2[2]), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[3]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC2_v2_3[0]), 
        .B(Red_MCInst_MC2_v1_3[0]), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC2_v0_3[0]), 
        .B(Red_MCInst_MC2_v3_3[0]), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[4]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC2_v2_3[1]), 
        .B(Red_MCInst_MC2_v1_3[1]), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC2_v0_3[1]), 
        .B(Red_MCInst_MC2_v3_3[1]), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[5]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC2_v2_3[2]), 
        .B(Red_MCInst_MC2_v1_3[2]), .ZN(Red_MCInst_MC2_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC2_v0_3[2]), 
        .B(Red_MCInst_MC2_v3_3[2]), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst_MC3_U3 ( .A(ShiftRowsOutput[16]), .Z(
        Red_MCInst_MC3_v2_1[1]) );
  BUF_X1 Red_MCInst_MC3_U2 ( .A(MCInst_MC3_v1_3[2]), .Z(Red_MCInst_MC3_v1_2[1]) );
  XOR2_X1 Red_MCInst_MC3_v0_2Inst_0_U1 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(Red_MCInst_MC3_v0_2[0]) );
  XOR2_X1 Red_MCInst_MC3_v0_3Inst_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_3[0]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U2 ( .A(Red_MCInst_MC3_v1_0Inst_0_n3), 
        .B(MCInst_MC3_v1_3[3]), .ZN(Red_MCInst_MC3_v1_0[0]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC3_v1_2Inst_0_U1 ( .A(Red_MCInst_MC3_v1_2[1]), .B(
        Red_MCInst_MC3_v1_1[2]), .Z(Red_MCInst_MC3_v1_2[0]) );
  XOR2_X1 Red_MCInst_MC3_v1_3Inst_0_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .Z(Red_MCInst_MC3_v1_3[0]) );
  XOR2_X1 Red_MCInst_MC3_v2_0Inst_0_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(Red_MCInst_MC3_v2_0[0]) );
  XOR2_X1 Red_MCInst_MC3_v2_1Inst_0_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_1[0]) );
  XNOR2_X1 Red_MCInst_MC3_v2_2Inst_0_U2 ( .A(Red_MCInst_MC3_v2_2Inst_0_n3), 
        .B(Red_MCInst_MC3_v2_2[1]), .ZN(Red_MCInst_MC3_v2_2[0]) );
  XNOR2_X1 Red_MCInst_MC3_v2_2Inst_0_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[2]), .ZN(Red_MCInst_MC3_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst_MC3_v2_3Inst_0_U2 ( .A(Red_MCInst_MC3_v2_3Inst_0_n3), 
        .B(Red_MCInst_MC3_v2_2[1]), .ZN(Red_MCInst_MC3_v2_3[0]) );
  XNOR2_X1 Red_MCInst_MC3_v2_3Inst_0_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[3]), .ZN(Red_MCInst_MC3_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst_MC3_v3_0Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_0[0]) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U3 ( .A(Red_MCInst_MC3_v3_2Inst_0_n6), 
        .B(Red_MCInst_MC3_v3_2Inst_0_n5), .ZN(Red_MCInst_MC3_v3_2[0]) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U2 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst_MC3_v3_3Inst_0_U1 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .Z(Red_MCInst_MC3_v3_3[0]) );
  XOR2_X1 Red_MCInst_MC3_v0_0Inst_1_U1 ( .A(Red_MCInst_MC3_v0_2[2]), .B(
        Red_MCInst_MC3_v0_1[0]), .Z(Red_MCInst_MC3_v0_0[1]) );
  XNOR2_X1 Red_MCInst_MC3_v0_1Inst_1_U2 ( .A(Red_MCInst_MC3_v0_1Inst_1_n3), 
        .B(Red_MCInst_MC3_v0_1[0]), .ZN(Red_MCInst_MC3_v0_1[1]) );
  XNOR2_X1 Red_MCInst_MC3_v0_1Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .ZN(Red_MCInst_MC3_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_2[1]) );
  XOR2_X1 Red_MCInst_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        MCInst_MC3_v0_3[3]), .Z(Red_MCInst_MC3_v0_3[1]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_1_U2 ( .A(Red_MCInst_MC3_v1_0Inst_1_n3), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_0[1]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_1Inst_1_U3 ( .A(Red_MCInst_MC3_v1_1Inst_1_n6), 
        .B(Red_MCInst_MC3_v1_1Inst_1_n5), .ZN(Red_MCInst_MC3_v1_1[1]) );
  XNOR2_X1 Red_MCInst_MC3_v1_1Inst_1_U2 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC3_v1_1Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .Z(Red_MCInst_MC3_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC3_v1_3Inst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[3]), .Z(Red_MCInst_MC3_v1_3[1]) );
  XOR2_X1 Red_MCInst_MC3_v2_0Inst_1_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_0[1]) );
  XOR2_X1 Red_MCInst_MC3_v2_3Inst_1_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(Red_MCInst_MC3_v2_3[1]) );
  XOR2_X1 Red_MCInst_MC3_v3_0Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .Z(Red_MCInst_MC3_v3_0[1]) );
  XNOR2_X1 Red_MCInst_MC3_v3_1Inst_1_U3 ( .A(Red_MCInst_MC3_v3_1Inst_1_n6), 
        .B(Red_MCInst_MC3_v3_1Inst_1_n5), .ZN(Red_MCInst_MC3_v3_1[1]) );
  XNOR2_X1 Red_MCInst_MC3_v3_1Inst_1_U2 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst_MC3_v3_1Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst_MC3_v3_2Inst_1_U1 ( .A(Red_MCInst_MC3_v3_3[2]), .B(
        MCInst_MC3_v3_0[3]), .Z(Red_MCInst_MC3_v3_2[1]) );
  XOR2_X1 Red_MCInst_MC3_v3_3Inst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_3[1]) );
  XNOR2_X1 Red_MCInst_MC3_v0_0Inst_2_U2 ( .A(Red_MCInst_MC3_v0_0Inst_2_n3), 
        .B(MCInst_MC3_v0_3[3]), .ZN(Red_MCInst_MC3_v0_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .ZN(Red_MCInst_MC3_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst_MC3_v0_1Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_1[2]) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_2_U3 ( .A(Red_MCInst_MC3_v0_3Inst_2_n6), 
        .B(Red_MCInst_MC3_v0_3Inst_2_n5), .ZN(Red_MCInst_MC3_v0_3[2]) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_2_U2 ( .A(MCInst_MC3_v0_3[3]), .B(
        Red_MCInst_MC3_v0_1[0]), .ZN(Red_MCInst_MC3_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v0_3Inst_2_U1 ( .A(Red_MCInst_MC3_v0_0[0]), .B(
        Red_MCInst_MC3_v0_2[2]), .Z(Red_MCInst_MC3_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_2_U2 ( .A(Red_MCInst_MC3_v1_0Inst_2_n3), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_2_U1 ( .A(Red_MCInst_MC3_v1_2[1]), .B(
        MCInst_MC3_v1_3[3]), .ZN(Red_MCInst_MC3_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_2Inst_2_U2 ( .A(Red_MCInst_MC3_v1_2Inst_2_n3), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_2[2]) );
  XNOR2_X1 Red_MCInst_MC3_v1_2Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_2_U3 ( .A(Red_MCInst_MC3_v1_3Inst_2_n6), 
        .B(Red_MCInst_MC3_v1_3Inst_2_n5), .ZN(Red_MCInst_MC3_v1_3[2]) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_2_U2 ( .A(MCInst_MC3_v1_3[3]), .B(
        Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v1_3Inst_2_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        Red_MCInst_MC3_v1_2[1]), .Z(Red_MCInst_MC3_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_2_U3 ( .A(Red_MCInst_MC3_v2_0Inst_2_n6), 
        .B(Red_MCInst_MC3_v2_0Inst_2_n5), .ZN(Red_MCInst_MC3_v2_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_2_U2 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .ZN(Red_MCInst_MC3_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v2_0Inst_2_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[2]), .Z(Red_MCInst_MC3_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst_MC3_v2_1Inst_2_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(Red_MCInst_MC3_v2_1[2]) );
  XOR2_X1 Red_MCInst_MC3_v2_2Inst_2_U1 ( .A(MCInst_MC3_v2_0[3]), .B(
        Red_MCInst_MC3_v2_2[1]), .Z(Red_MCInst_MC3_v2_2[2]) );
  XOR2_X1 Red_MCInst_MC3_v2_3Inst_2_U1 ( .A(Red_MCInst_MC3_v2_1[1]), .B(
        MCInst_MC3_v2_0[3]), .Z(Red_MCInst_MC3_v2_3[2]) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_2_U3 ( .A(Red_MCInst_MC3_v3_0Inst_2_n6), 
        .B(Red_MCInst_MC3_v3_0Inst_2_n5), .ZN(Red_MCInst_MC3_v3_0[2]) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_2_U2 ( .A(MCInst_MC3_v3_0[3]), .B(
        Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst_MC3_v3_0Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_2_U2 ( .A(Red_MCInst_MC3_v3_2Inst_2_n3), 
        .B(Red_MCInst_MC3_v3_1[2]), .ZN(Red_MCInst_MC3_v3_2[2]) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_2_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        MCInst_MC3_v3_0[3]), .ZN(Red_MCInst_MC3_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output[36]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_0[0]), 
        .B(Red_MCInst_MC3_v1_0[0]), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), 
        .B(Red_MCInst_MC3_v3_0[0]), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output[37]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_0[1]), 
        .B(Red_MCInst_MC3_v1_0[1]), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_0[1]), 
        .B(Red_MCInst_MC3_v3_0[1]), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output[38]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_0[2]), 
        .B(Red_MCInst_MC3_v1_0[2]), .ZN(Red_MCInst_MC3_r0Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_0[2]), 
        .B(Red_MCInst_MC3_v3_0[2]), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output[24]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_1[0]), 
        .B(Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_1[0]), 
        .B(Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output[25]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_1[1]), 
        .B(Red_MCInst_MC3_v1_1[1]), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_1[1]), 
        .B(Red_MCInst_MC3_v3_1[1]), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output[26]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_1[2]), 
        .B(Red_MCInst_MC3_v1_1[2]), .ZN(Red_MCInst_MC3_r1Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_1[2]), 
        .B(Red_MCInst_MC3_v3_1[2]), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output[12]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_2[0]), 
        .B(Red_MCInst_MC3_v1_2[0]), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_2[0]), 
        .B(Red_MCInst_MC3_v3_2[0]), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output[13]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_2[1]), 
        .B(Red_MCInst_MC3_v1_2[1]), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_2[1]), 
        .B(Red_MCInst_MC3_v3_2[1]), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output[14]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_2[2]), 
        .B(Red_MCInst_MC3_v1_2[2]), .ZN(Red_MCInst_MC3_r2Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), 
        .B(Red_MCInst_MC3_v3_2[2]), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output[0]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst_MC3_v2_3[0]), 
        .B(Red_MCInst_MC3_v1_3[0]), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_0_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst_MC3_v0_3[0]), 
        .B(Red_MCInst_MC3_v3_3[0]), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output[1]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst_MC3_v2_3[1]), 
        .B(Red_MCInst_MC3_v1_3[1]), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_1_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst_MC3_v0_3[1]), 
        .B(Red_MCInst_MC3_v3_3[1]), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output[2]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst_MC3_v2_3[2]), 
        .B(Red_MCInst_MC3_v1_3[2]), .ZN(Red_MCInst_MC3_r3Inst_XORInst_0_2_n7)
         );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst_MC3_v0_3[2]), 
        .B(Red_MCInst_MC3_v3_3[2]), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_2_n8)
         );
  DFF_X1 RedStateReg_s_current_state_reg_0_ ( .D(Red_MC_output[0]), .CK(clk), 
        .Q(Red_SubCellInput2[0]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_1_ ( .D(Red_MC_output[1]), .CK(clk), 
        .Q(Red_SubCellInput2[1]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_2_ ( .D(Red_MC_output[2]), .CK(clk), 
        .Q(Red_SubCellInput2[2]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_3_ ( .D(Red_MC_output[3]), .CK(clk), 
        .Q(Red_SubCellInput2[3]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_4_ ( .D(Red_MC_output[4]), .CK(clk), 
        .Q(Red_SubCellInput2[4]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_5_ ( .D(Red_MC_output[5]), .CK(clk), 
        .Q(Red_SubCellInput2[5]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_6_ ( .D(Red_MC_output[6]), .CK(clk), 
        .Q(Red_SubCellInput2[6]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_7_ ( .D(Red_MC_output[7]), .CK(clk), 
        .Q(Red_SubCellInput2[7]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_8_ ( .D(Red_MC_output[8]), .CK(clk), 
        .Q(Red_SubCellInput2[8]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_9_ ( .D(Red_MC_output[9]), .CK(clk), 
        .Q(Red_SubCellInput2[9]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_10_ ( .D(Red_MC_output[10]), .CK(clk), 
        .Q(Red_SubCellInput2[10]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_11_ ( .D(Red_MC_output[11]), .CK(clk), 
        .Q(Red_SubCellInput2[11]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_12_ ( .D(Red_MC_output[12]), .CK(clk), 
        .Q(Red_SubCellInput2[12]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_13_ ( .D(Red_MC_output[13]), .CK(clk), 
        .Q(Red_SubCellInput2[13]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_14_ ( .D(Red_MC_output[14]), .CK(clk), 
        .Q(Red_SubCellInput2[14]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_15_ ( .D(Red_MC_output[15]), .CK(clk), 
        .Q(Red_SubCellInput2[15]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_16_ ( .D(Red_MC_output[16]), .CK(clk), 
        .Q(Red_SubCellInput2[16]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_17_ ( .D(Red_MC_output[17]), .CK(clk), 
        .Q(Red_SubCellInput2[17]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_18_ ( .D(Red_MC_output[18]), .CK(clk), 
        .Q(Red_SubCellInput2[18]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_19_ ( .D(Red_MC_output[19]), .CK(clk), 
        .Q(Red_SubCellInput2[19]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_20_ ( .D(Red_MC_output[20]), .CK(clk), 
        .Q(Red_SubCellInput2[20]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_21_ ( .D(Red_MC_output[21]), .CK(clk), 
        .Q(Red_SubCellInput2[21]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_22_ ( .D(Red_MC_output[22]), .CK(clk), 
        .Q(Red_SubCellInput2[22]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_23_ ( .D(Red_MC_output[23]), .CK(clk), 
        .Q(Red_SubCellInput2[23]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_24_ ( .D(Red_MC_output[24]), .CK(clk), 
        .Q(Red_SubCellInput2[24]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_25_ ( .D(Red_MC_output[25]), .CK(clk), 
        .Q(Red_SubCellInput2[25]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_26_ ( .D(Red_MC_output[26]), .CK(clk), 
        .Q(Red_SubCellInput2[26]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_27_ ( .D(Red_MC_output[27]), .CK(clk), 
        .Q(Red_SubCellInput2[27]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_28_ ( .D(Red_MC_output[28]), .CK(clk), 
        .Q(Red_SubCellInput2[28]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_29_ ( .D(Red_MC_output[29]), .CK(clk), 
        .Q(Red_SubCellInput2[29]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_30_ ( .D(Red_MC_output[30]), .CK(clk), 
        .Q(Red_SubCellInput2[30]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_31_ ( .D(Red_MC_output[31]), .CK(clk), 
        .Q(Red_SubCellInput2[31]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_32_ ( .D(Red_MC_output[32]), .CK(clk), 
        .Q(Red_SubCellInput2[32]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_33_ ( .D(Red_MC_output[33]), .CK(clk), 
        .Q(Red_SubCellInput2[33]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_34_ ( .D(Red_MC_output[34]), .CK(clk), 
        .Q(Red_SubCellInput2[34]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_35_ ( .D(Red_MC_output[35]), .CK(clk), 
        .Q(Red_SubCellInput2[35]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_36_ ( .D(Red_MC_output[36]), .CK(clk), 
        .Q(Red_SubCellInput2[36]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_37_ ( .D(Red_MC_output[37]), .CK(clk), 
        .Q(Red_SubCellInput2[37]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_38_ ( .D(Red_MC_output[38]), .CK(clk), 
        .Q(Red_SubCellInput2[38]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_39_ ( .D(Red_MC_output[39]), .CK(clk), 
        .Q(Red_SubCellInput2[39]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_40_ ( .D(Red_MC_output[40]), .CK(clk), 
        .Q(Red_SubCellInput2[40]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_41_ ( .D(Red_MC_output[41]), .CK(clk), 
        .Q(Red_SubCellInput2[41]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_42_ ( .D(Red_MC_output[42]), .CK(clk), 
        .Q(Red_SubCellInput2[42]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_43_ ( .D(Red_MC_output[43]), .CK(clk), 
        .Q(Red_SubCellInput2[43]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_44_ ( .D(Red_MC_output[44]), .CK(clk), 
        .Q(Red_SubCellInput2[44]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_45_ ( .D(Red_MC_output[45]), .CK(clk), 
        .Q(Red_SubCellInput2[45]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_46_ ( .D(Red_MC_output[46]), .CK(clk), 
        .Q(Red_SubCellInput2[46]), .QN() );
  DFF_X1 RedStateReg_s_current_state_reg_47_ ( .D(Red_MC_output[47]), .CK(clk), 
        .Q(Red_SubCellInput2[47]), .QN() );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[9])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U4 ( .A1(SubCellInput2[2]), .A2(
        SubCellInput2[3]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U3 ( .A1(SubCellInput2[0]), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U2 ( .A1(SubCellInput2[2]), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U1 ( .A(SubCellInput2[1]), .B(
        SubCellInput2[3]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[10])
         );
  OR2_X1 Red_SubCellInst2_LFInst_0_LFInst_1_U2 ( .A1(SubCellInput2[3]), .A2(
        SubCellInput2[2]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_1_U1 ( .A1(SubCellInput2[1]), .A2(
        SubCellInput2[3]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[11])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_2_n15), .A2(SubCellInput2[3]), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_2_n14), .A2(SubCellInput2[2]), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U4 ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U2 ( .A(SubCellInput2[1]), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_0_LFInst_2_U1 ( .A(SubCellInput2[0]), .B(
        SubCellInput2[2]), .Z(Red_SubCellInst2_LFInst_0_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[0])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U4 ( .A1(SubCellInput2[6]), .A2(
        SubCellInput2[7]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U3 ( .A1(SubCellInput2[4]), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U2 ( .A1(SubCellInput2[6]), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U1 ( .A(SubCellInput2[5]), .B(
        SubCellInput2[7]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[1])
         );
  OR2_X1 Red_SubCellInst2_LFInst_1_LFInst_1_U2 ( .A1(SubCellInput2[7]), .A2(
        SubCellInput2[6]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_1_U1 ( .A1(SubCellInput2[5]), .A2(
        SubCellInput2[7]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_2_n14), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_2_n13), .ZN(Red_ShiftRowsOutput2[2])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_2_n12), .A2(SubCellInput2[7]), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_2_n11), .A2(SubCellInput2[6]), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U4 ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_2_n11) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_2_n10), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_2_n9), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_2_n14) );
  INV_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U2 ( .A(SubCellInput2[5]), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_2_n9) );
  XOR2_X1 Red_SubCellInst2_LFInst_1_LFInst_2_U1 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[6]), .Z(Red_SubCellInst2_LFInst_1_LFInst_2_n10) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[3])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U4 ( .A1(SubCellInput2[10]), 
        .A2(SubCellInput2[11]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U3 ( .A1(SubCellInput2[8]), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U2 ( .A1(SubCellInput2[10]), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U1 ( .A(SubCellInput2[9]), .B(
        SubCellInput2[11]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[4])
         );
  OR2_X1 Red_SubCellInst2_LFInst_2_LFInst_1_U2 ( .A1(SubCellInput2[11]), .A2(
        SubCellInput2[10]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_1_U1 ( .A1(SubCellInput2[9]), .A2(
        SubCellInput2[11]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[5])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_2_n15), .A2(SubCellInput2[11]), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_2_n14), .A2(SubCellInput2[10]), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U4 ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U2 ( .A(SubCellInput2[9]), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_2_LFInst_2_U1 ( .A(SubCellInput2[8]), .B(
        SubCellInput2[10]), .Z(Red_SubCellInst2_LFInst_2_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[6])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U4 ( .A1(SubCellInput2[14]), 
        .A2(SubCellInput2[15]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U3 ( .A1(SubCellInput2[12]), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U2 ( .A1(SubCellInput2[14]), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U1 ( .A(SubCellInput2[13]), .B(
        SubCellInput2[15]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[7])
         );
  OR2_X1 Red_SubCellInst2_LFInst_3_LFInst_1_U2 ( .A1(SubCellInput2[15]), .A2(
        SubCellInput2[14]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_1_U1 ( .A1(SubCellInput2[13]), 
        .A2(SubCellInput2[15]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[8])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_2_n15), .A2(SubCellInput2[15]), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_2_n14), .A2(SubCellInput2[14]), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U4 ( .A1(SubCellInput2[12]), 
        .A2(SubCellInput2[13]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U2 ( .A(SubCellInput2[13]), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_3_LFInst_2_U1 ( .A(SubCellInput2[12]), .B(
        SubCellInput2[14]), .Z(Red_SubCellInst2_LFInst_3_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[18])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U4 ( .A1(SubCellInput2[18]), 
        .A2(SubCellInput2[19]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U3 ( .A1(SubCellInput2[16]), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U2 ( .A1(SubCellInput2[18]), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U1 ( .A(SubCellInput2[17]), .B(
        SubCellInput2[19]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[19])
         );
  OR2_X1 Red_SubCellInst2_LFInst_4_LFInst_1_U2 ( .A1(SubCellInput2[19]), .A2(
        SubCellInput2[18]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_1_U1 ( .A1(SubCellInput2[17]), 
        .A2(SubCellInput2[19]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_2_n14), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[20])
         );
  OR2_X1 Red_SubCellInst2_LFInst_4_LFInst_2_U5 ( .A1(SubCellInput2[17]), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_2_n15), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst2_LFInst_4_LFInst_2_U4 ( .A(SubCellInput2[18]), .B(
        SubCellInput2[16]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_2_n13), .A2(SubCellInput2[19]), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_2_U2 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_2_n12), .A2(SubCellInput2[18]), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_2_U1 ( .A1(SubCellInput2[16]), 
        .A2(SubCellInput2[17]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[21])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U4 ( .A1(SubCellInput2[22]), 
        .A2(SubCellInput2[23]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U3 ( .A1(SubCellInput2[20]), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U2 ( .A1(SubCellInput2[22]), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U1 ( .A(SubCellInput2[21]), .B(
        SubCellInput2[23]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[22])
         );
  OR2_X1 Red_SubCellInst2_LFInst_5_LFInst_1_U2 ( .A1(SubCellInput2[23]), .A2(
        SubCellInput2[22]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_1_U1 ( .A1(SubCellInput2[21]), 
        .A2(SubCellInput2[23]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[23])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_2_n15), .A2(SubCellInput2[23]), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_2_n14), .A2(SubCellInput2[22]), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U4 ( .A1(SubCellInput2[20]), 
        .A2(SubCellInput2[21]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U2 ( .A(SubCellInput2[21]), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_5_LFInst_2_U1 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[22]), .Z(Red_SubCellInst2_LFInst_5_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[12])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U4 ( .A1(SubCellInput2[26]), 
        .A2(SubCellInput2[27]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U3 ( .A1(SubCellInput2[24]), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U2 ( .A1(SubCellInput2[26]), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U1 ( .A(SubCellInput2[25]), .B(
        SubCellInput2[27]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[13])
         );
  OR2_X1 Red_SubCellInst2_LFInst_6_LFInst_1_U2 ( .A1(SubCellInput2[27]), .A2(
        SubCellInput2[26]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_1_U1 ( .A1(SubCellInput2[25]), 
        .A2(SubCellInput2[27]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[14])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_2_n15), .A2(SubCellInput2[27]), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_2_n14), .A2(SubCellInput2[26]), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U4 ( .A1(SubCellInput2[24]), 
        .A2(SubCellInput2[25]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U2 ( .A(SubCellInput2[25]), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_6_LFInst_2_U1 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[26]), .Z(Red_SubCellInst2_LFInst_6_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[15])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U4 ( .A1(SubCellInput2[30]), 
        .A2(SubCellInput2[31]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U3 ( .A1(SubCellInput2[28]), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U2 ( .A1(SubCellInput2[30]), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U1 ( .A(SubCellInput2[29]), .B(
        SubCellInput2[31]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[16])
         );
  OR2_X1 Red_SubCellInst2_LFInst_7_LFInst_1_U2 ( .A1(SubCellInput2[31]), .A2(
        SubCellInput2[30]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_1_U1 ( .A1(SubCellInput2[29]), 
        .A2(SubCellInput2[31]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[17])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_2_n15), .A2(SubCellInput2[31]), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_2_n14), .A2(SubCellInput2[30]), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U4 ( .A1(SubCellInput2[28]), 
        .A2(SubCellInput2[29]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U2 ( .A(SubCellInput2[29]), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_7_LFInst_2_U1 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[30]), .Z(Red_SubCellInst2_LFInst_7_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[27])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U4 ( .A1(SubCellInput2[34]), 
        .A2(SubCellInput2[35]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U3 ( .A1(SubCellInput2[32]), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U2 ( .A1(SubCellInput2[34]), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U1 ( .A(SubCellInput2[33]), .B(
        SubCellInput2[35]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[28])
         );
  OR2_X1 Red_SubCellInst2_LFInst_8_LFInst_1_U2 ( .A1(SubCellInput2[35]), .A2(
        SubCellInput2[34]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_1_U1 ( .A1(SubCellInput2[33]), 
        .A2(SubCellInput2[35]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_2_n14), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_2_n13), .ZN(Red_ShiftRowsOutput2[29])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_2_n12), .A2(SubCellInput2[35]), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_2_n11), .A2(SubCellInput2[34]), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U4 ( .A1(SubCellInput2[32]), 
        .A2(SubCellInput2[33]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_2_n11) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_2_n10), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_2_n9), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_2_n14) );
  INV_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U2 ( .A(SubCellInput2[33]), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_2_n9) );
  XOR2_X1 Red_SubCellInst2_LFInst_8_LFInst_2_U1 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[34]), .Z(Red_SubCellInst2_LFInst_8_LFInst_2_n10) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[30])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U4 ( .A1(SubCellInput2[38]), 
        .A2(SubCellInput2[39]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n11) );
  OR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U3 ( .A1(SubCellInput2[36]), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U2 ( .A1(SubCellInput2[38]), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U1 ( .A(SubCellInput2[37]), .B(
        SubCellInput2[39]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[31])
         );
  OR2_X1 Red_SubCellInst2_LFInst_9_LFInst_1_U2 ( .A1(SubCellInput2[39]), .A2(
        SubCellInput2[38]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_1_U1 ( .A1(SubCellInput2[37]), 
        .A2(SubCellInput2[39]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_2_n14), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[32])
         );
  OR2_X1 Red_SubCellInst2_LFInst_9_LFInst_2_U5 ( .A1(SubCellInput2[37]), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_2_n15), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst2_LFInst_9_LFInst_2_U4 ( .A(SubCellInput2[38]), .B(
        SubCellInput2[36]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_2_n13), .A2(SubCellInput2[39]), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_2_U2 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_2_n12), .A2(SubCellInput2[38]), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_2_U1 ( .A1(SubCellInput2[36]), 
        .A2(SubCellInput2[37]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[33]) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U4 ( .A1(SubCellInput2[42]), 
        .A2(SubCellInput2[43]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U3 ( .A1(SubCellInput2[40]), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U2 ( .A1(SubCellInput2[42]), 
        .A2(Red_SubCellInst2_LFInst_10_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U1 ( .A(SubCellInput2[41]), .B(
        SubCellInput2[43]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[34])
         );
  OR2_X1 Red_SubCellInst2_LFInst_10_LFInst_1_U2 ( .A1(SubCellInput2[43]), .A2(
        SubCellInput2[42]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_1_U1 ( .A1(SubCellInput2[41]), 
        .A2(SubCellInput2[43]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[35]) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_2_n15), .A2(SubCellInput2[43]), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_2_n14), .A2(SubCellInput2[42]), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U4 ( .A1(SubCellInput2[40]), 
        .A2(SubCellInput2[41]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U2 ( .A(SubCellInput2[41]), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_10_LFInst_2_U1 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[42]), .Z(Red_SubCellInst2_LFInst_10_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[24]) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U4 ( .A1(SubCellInput2[46]), 
        .A2(SubCellInput2[47]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U3 ( .A1(SubCellInput2[44]), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U2 ( .A1(SubCellInput2[46]), 
        .A2(Red_SubCellInst2_LFInst_11_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U1 ( .A(SubCellInput2[45]), .B(
        SubCellInput2[47]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[25])
         );
  OR2_X1 Red_SubCellInst2_LFInst_11_LFInst_1_U2 ( .A1(SubCellInput2[47]), .A2(
        SubCellInput2[46]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_1_U1 ( .A1(SubCellInput2[45]), 
        .A2(SubCellInput2[47]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[26]) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_2_n15), .A2(SubCellInput2[47]), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_2_n14), .A2(SubCellInput2[46]), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U4 ( .A1(SubCellInput2[44]), 
        .A2(SubCellInput2[45]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U2 ( .A(SubCellInput2[45]), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_11_LFInst_2_U1 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[46]), .Z(Red_SubCellInst2_LFInst_11_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[36]) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U4 ( .A1(SubCellInput2[50]), 
        .A2(SubCellInput2[51]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U3 ( .A1(SubCellInput2[48]), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U2 ( .A1(SubCellInput2[50]), 
        .A2(Red_SubCellInst2_LFInst_12_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U1 ( .A(SubCellInput2[49]), .B(
        SubCellInput2[51]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[37])
         );
  OR2_X1 Red_SubCellInst2_LFInst_12_LFInst_1_U2 ( .A1(SubCellInput2[51]), .A2(
        SubCellInput2[50]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_1_U1 ( .A1(SubCellInput2[49]), 
        .A2(SubCellInput2[51]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_2_n16), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_2_n15), .ZN(Red_ShiftRowsOutput2[38]) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_2_n14), .A2(SubCellInput2[51]), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_2_U4 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_2_n13), .A2(SubCellInput2[50]), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_2_U3 ( .A1(SubCellInput2[48]), 
        .A2(SubCellInput2[49]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_2_n13)
         );
  OR2_X1 Red_SubCellInst2_LFInst_12_LFInst_2_U2 ( .A1(SubCellInput2[49]), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst2_LFInst_12_LFInst_2_U1 ( .A(SubCellInput2[50]), .B(
        SubCellInput2[48]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[39]) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U4 ( .A1(SubCellInput2[54]), 
        .A2(SubCellInput2[55]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U3 ( .A1(SubCellInput2[52]), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U2 ( .A1(SubCellInput2[54]), 
        .A2(Red_SubCellInst2_LFInst_13_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U1 ( .A(SubCellInput2[53]), .B(
        SubCellInput2[55]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[40])
         );
  OR2_X1 Red_SubCellInst2_LFInst_13_LFInst_1_U2 ( .A1(SubCellInput2[55]), .A2(
        SubCellInput2[54]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_1_U1 ( .A1(SubCellInput2[53]), 
        .A2(SubCellInput2[55]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[41]) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_2_n15), .A2(SubCellInput2[55]), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_2_n14), .A2(SubCellInput2[54]), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U4 ( .A1(SubCellInput2[52]), 
        .A2(SubCellInput2[53]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U2 ( .A(SubCellInput2[53]), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_13_LFInst_2_U1 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[54]), .Z(Red_SubCellInst2_LFInst_13_LFInst_2_n13) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[42]) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U4 ( .A1(SubCellInput2[58]), 
        .A2(SubCellInput2[59]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U3 ( .A1(SubCellInput2[56]), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U2 ( .A1(SubCellInput2[58]), 
        .A2(Red_SubCellInst2_LFInst_14_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U1 ( .A(SubCellInput2[57]), .B(
        SubCellInput2[59]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[43])
         );
  OR2_X1 Red_SubCellInst2_LFInst_14_LFInst_1_U2 ( .A1(SubCellInput2[59]), .A2(
        SubCellInput2[58]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_1_U1 ( .A1(SubCellInput2[57]), 
        .A2(SubCellInput2[59]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_2_n16), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_2_n15), .ZN(Red_ShiftRowsOutput2[44]) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_2_n14), .A2(SubCellInput2[59]), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_2_U4 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_2_n13), .A2(SubCellInput2[58]), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_2_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_2_U3 ( .A1(SubCellInput2[56]), 
        .A2(SubCellInput2[57]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_2_n13)
         );
  OR2_X1 Red_SubCellInst2_LFInst_14_LFInst_2_U2 ( .A1(SubCellInput2[57]), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_2_n16) );
  XNOR2_X1 Red_SubCellInst2_LFInst_14_LFInst_2_U1 ( .A(SubCellInput2[58]), .B(
        SubCellInput2[56]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_2_n12) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_0_n12), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_0_n11), .ZN(Red_ShiftRowsOutput2[45]) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U4 ( .A1(SubCellInput2[62]), 
        .A2(SubCellInput2[63]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n11)
         );
  OR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U3 ( .A1(SubCellInput2[60]), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_0_n10), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n12) );
  NOR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U2 ( .A1(SubCellInput2[62]), 
        .A2(Red_SubCellInst2_LFInst_15_LFInst_0_n9), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n10) );
  XNOR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U1 ( .A(SubCellInput2[61]), .B(
        SubCellInput2[63]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n9) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_1_U3 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_1_n6), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_1_n5), .ZN(Red_ShiftRowsOutput2[46])
         );
  OR2_X1 Red_SubCellInst2_LFInst_15_LFInst_1_U2 ( .A1(SubCellInput2[63]), .A2(
        SubCellInput2[62]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_1_n5) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_1_U1 ( .A1(SubCellInput2[61]), 
        .A2(SubCellInput2[63]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_1_n6) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U7 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_2_n17), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_2_n16), .ZN(Red_ShiftRowsOutput2[47]) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U6 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_2_n15), .A2(SubCellInput2[63]), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_2_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U5 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_2_n14), .A2(SubCellInput2[62]), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_2_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U4 ( .A1(SubCellInput2[60]), 
        .A2(SubCellInput2[61]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_2_n14)
         );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U3 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_2_n13), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_2_n12), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_2_n17) );
  INV_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U2 ( .A(SubCellInput2[61]), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_2_n12) );
  XOR2_X1 Red_SubCellInst2_LFInst_15_LFInst_2_U1 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[62]), .Z(Red_SubCellInst2_LFInst_15_LFInst_2_n13) );
  BUF_X1 Red_MCInst2_MC0_U3 ( .A(ShiftRowsOutput2[28]), .Z(
        Red_MCInst2_MC0_v2_1[1]) );
  BUF_X1 Red_MCInst2_MC0_U2 ( .A(MCInst2_MC0_v1_3[2]), .Z(
        Red_MCInst2_MC0_v1_2[1]) );
  XOR2_X1 Red_MCInst2_MC0_v0_2Inst_0_U1 ( .A(MCInst2_MC0_v0_3[3]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(Red_MCInst2_MC0_v0_2[0]) );
  XOR2_X1 Red_MCInst2_MC0_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_2[2]), .Z(Red_MCInst2_MC0_v0_3[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC0_v1_0Inst_0_n3), 
        .B(MCInst2_MC0_v1_3[3]), .ZN(Red_MCInst2_MC0_v1_0[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_2[1]), .ZN(Red_MCInst2_MC0_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC0_v1_2Inst_0_U1 ( .A(Red_MCInst2_MC0_v1_2[1]), .B(
        Red_MCInst2_MC0_v1_1[2]), .Z(Red_MCInst2_MC0_v1_2[0]) );
  XOR2_X1 Red_MCInst2_MC0_v1_3Inst_0_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_2[1]), .Z(Red_MCInst2_MC0_v1_3[0]) );
  XOR2_X1 Red_MCInst2_MC0_v2_0Inst_0_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(Red_MCInst2_MC0_v2_0[0]) );
  XOR2_X1 Red_MCInst2_MC0_v2_1Inst_0_U1 ( .A(MCInst2_MC0_v2_0[2]), .B(
        MCInst2_MC0_v2_0[3]), .Z(Red_MCInst2_MC0_v2_1[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v2_2Inst_0_U2 ( .A(Red_MCInst2_MC0_v2_2Inst_0_n3), 
        .B(Red_MCInst2_MC0_v2_2[1]), .ZN(Red_MCInst2_MC0_v2_2[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v2_2Inst_0_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v2_0[2]), .ZN(Red_MCInst2_MC0_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v2_3Inst_0_U2 ( .A(Red_MCInst2_MC0_v2_3Inst_0_n3), 
        .B(Red_MCInst2_MC0_v2_2[1]), .ZN(Red_MCInst2_MC0_v2_3[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v2_3Inst_0_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v2_0[3]), .ZN(Red_MCInst2_MC0_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC0_v3_0Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_v3_0[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U3 ( .A(Red_MCInst2_MC0_v3_2Inst_0_n6), 
        .B(Red_MCInst2_MC0_v3_2Inst_0_n5), .ZN(Red_MCInst2_MC0_v3_2[0]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U2 ( .A(MCInst2_MC0_v3_0[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .ZN(Red_MCInst2_MC0_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC0_v3_3Inst_0_U1 ( .A(MCInst2_MC0_v3_0[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .Z(Red_MCInst2_MC0_v3_3[0]) );
  XOR2_X1 Red_MCInst2_MC0_v0_0Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), .B(
        Red_MCInst2_MC0_v0_1[0]), .Z(Red_MCInst2_MC0_v0_0[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v0_1Inst_1_U2 ( .A(Red_MCInst2_MC0_v0_1Inst_1_n3), 
        .B(Red_MCInst2_MC0_v0_1[0]), .ZN(Red_MCInst2_MC0_v0_1[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        MCInst2_MC0_v0_3[3]), .ZN(Red_MCInst2_MC0_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst2_MC0_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_2[2]), .Z(Red_MCInst2_MC0_v0_2[1]) );
  XOR2_X1 Red_MCInst2_MC0_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        MCInst2_MC0_v0_3[3]), .Z(Red_MCInst2_MC0_v0_3[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_1_U2 ( .A(Red_MCInst2_MC0_v1_0Inst_1_n3), 
        .B(Red_MCInst2_MC0_v1_1[2]), .ZN(Red_MCInst2_MC0_v1_0[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_2[1]), .ZN(Red_MCInst2_MC0_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v1_1Inst_1_U3 ( .A(Red_MCInst2_MC0_v1_1Inst_1_n6), 
        .B(Red_MCInst2_MC0_v1_1Inst_1_n5), .ZN(Red_MCInst2_MC0_v1_1[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_1Inst_1_U2 ( .A(MCInst2_MC0_v1_3[3]), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(Red_MCInst2_MC0_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC0_v1_1Inst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_2[1]), .Z(Red_MCInst2_MC0_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC0_v1_3Inst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        MCInst2_MC0_v1_3[3]), .Z(Red_MCInst2_MC0_v1_3[1]) );
  XOR2_X1 Red_MCInst2_MC0_v2_0Inst_1_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v2_0[3]), .Z(Red_MCInst2_MC0_v2_0[1]) );
  XOR2_X1 Red_MCInst2_MC0_v2_3Inst_1_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        Red_MCInst2_MC0_v2_2[1]), .Z(Red_MCInst2_MC0_v2_3[1]) );
  XOR2_X1 Red_MCInst2_MC0_v3_0Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[3]), .Z(Red_MCInst2_MC0_v3_0[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_1Inst_1_U3 ( .A(Red_MCInst2_MC0_v3_1Inst_1_n6), 
        .B(Red_MCInst2_MC0_v3_1Inst_1_n5), .ZN(Red_MCInst2_MC0_v3_1[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_1Inst_1_U2 ( .A(MCInst2_MC0_v3_0[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .ZN(Red_MCInst2_MC0_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC0_v3_1Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC0_v3_2Inst_1_U1 ( .A(Red_MCInst2_MC0_v3_3[2]), .B(
        MCInst2_MC0_v3_0[3]), .Z(Red_MCInst2_MC0_v3_2[1]) );
  XOR2_X1 Red_MCInst2_MC0_v3_3Inst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_v3_3[1]) );
  XNOR2_X1 Red_MCInst2_MC0_v0_0Inst_2_U2 ( .A(Red_MCInst2_MC0_v0_0Inst_2_n3), 
        .B(MCInst2_MC0_v0_3[3]), .ZN(Red_MCInst2_MC0_v0_0[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_2[2]), .ZN(Red_MCInst2_MC0_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst2_MC0_v0_1Inst_2_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_2[2]), .Z(Red_MCInst2_MC0_v0_1[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v0_3Inst_2_U3 ( .A(Red_MCInst2_MC0_v0_3Inst_2_n6), 
        .B(Red_MCInst2_MC0_v0_3Inst_2_n5), .ZN(Red_MCInst2_MC0_v0_3[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v0_3Inst_2_U2 ( .A(MCInst2_MC0_v0_3[3]), .B(
        Red_MCInst2_MC0_v0_1[0]), .ZN(Red_MCInst2_MC0_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC0_v0_3Inst_2_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), .B(
        Red_MCInst2_MC0_v0_2[2]), .Z(Red_MCInst2_MC0_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_2_U2 ( .A(Red_MCInst2_MC0_v1_0Inst_2_n3), 
        .B(Red_MCInst2_MC0_v1_1[2]), .ZN(Red_MCInst2_MC0_v1_0[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_2_U1 ( .A(Red_MCInst2_MC0_v1_2[1]), .B(
        MCInst2_MC0_v1_3[3]), .ZN(Red_MCInst2_MC0_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v1_2Inst_2_U2 ( .A(Red_MCInst2_MC0_v1_2Inst_2_n3), 
        .B(Red_MCInst2_MC0_v1_1[2]), .ZN(Red_MCInst2_MC0_v1_2[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_2Inst_2_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_2[1]), .ZN(Red_MCInst2_MC0_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC0_v1_3Inst_2_U3 ( .A(Red_MCInst2_MC0_v1_3Inst_2_n6), 
        .B(Red_MCInst2_MC0_v1_3Inst_2_n5), .ZN(Red_MCInst2_MC0_v1_3[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v1_3Inst_2_U2 ( .A(MCInst2_MC0_v1_3[3]), .B(
        Red_MCInst2_MC0_v1_1[2]), .ZN(Red_MCInst2_MC0_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC0_v1_3Inst_2_U1 ( .A(MCInst2_MC0_v1_0_0_), .B(
        Red_MCInst2_MC0_v1_2[1]), .Z(Red_MCInst2_MC0_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC0_v2_0Inst_2_U3 ( .A(Red_MCInst2_MC0_v2_0Inst_2_n6), 
        .B(Red_MCInst2_MC0_v2_0Inst_2_n5), .ZN(Red_MCInst2_MC0_v2_0[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v2_0Inst_2_U2 ( .A(MCInst2_MC0_v2_0[3]), .B(
        Red_MCInst2_MC0_v2_2[1]), .ZN(Red_MCInst2_MC0_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC0_v2_0Inst_2_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v2_0[2]), .Z(Red_MCInst2_MC0_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst2_MC0_v2_1Inst_2_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        Red_MCInst2_MC0_v2_2[1]), .Z(Red_MCInst2_MC0_v2_1[2]) );
  XOR2_X1 Red_MCInst2_MC0_v2_2Inst_2_U1 ( .A(MCInst2_MC0_v2_0[3]), .B(
        Red_MCInst2_MC0_v2_2[1]), .Z(Red_MCInst2_MC0_v2_2[2]) );
  XOR2_X1 Red_MCInst2_MC0_v2_3Inst_2_U1 ( .A(Red_MCInst2_MC0_v2_1[1]), .B(
        MCInst2_MC0_v2_0[3]), .Z(Red_MCInst2_MC0_v2_3[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_0Inst_2_U3 ( .A(Red_MCInst2_MC0_v3_0Inst_2_n6), 
        .B(Red_MCInst2_MC0_v3_0Inst_2_n5), .ZN(Red_MCInst2_MC0_v3_0[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_0Inst_2_U2 ( .A(MCInst2_MC0_v3_0[3]), .B(
        Red_MCInst2_MC0_v3_1[2]), .ZN(Red_MCInst2_MC0_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC0_v3_0Inst_2_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_2_U2 ( .A(Red_MCInst2_MC0_v3_2Inst_2_n3), 
        .B(Red_MCInst2_MC0_v3_1[2]), .ZN(Red_MCInst2_MC0_v3_2[2]) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_2_U1 ( .A(MCInst2_MC0_v3_2[3]), .B(
        MCInst2_MC0_v3_0[3]), .ZN(Red_MCInst2_MC0_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[45]) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_0[0]), 
        .B(Red_MCInst2_MC0_v1_0[0]), .ZN(Red_MCInst2_MC0_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), 
        .B(Red_MCInst2_MC0_v3_0[0]), .Z(Red_MCInst2_MC0_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC0_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC0_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[46]) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC0_v2_0[1]), 
        .B(Red_MCInst2_MC0_v1_0[1]), .ZN(Red_MCInst2_MC0_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC0_v0_0[1]), 
        .B(Red_MCInst2_MC0_v3_0[1]), .Z(Red_MCInst2_MC0_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC0_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC0_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[47]) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC0_v2_0[2]), 
        .B(Red_MCInst2_MC0_v1_0[2]), .ZN(Red_MCInst2_MC0_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC0_v0_0[2]), 
        .B(Red_MCInst2_MC0_v3_0[2]), .Z(Red_MCInst2_MC0_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[33]) );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_1[0]), 
        .B(Red_MCInst2_MC0_v1_2[1]), .ZN(Red_MCInst2_MC0_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_1[0]), 
        .B(Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC0_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC0_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[34]) );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC0_v2_1[1]), 
        .B(Red_MCInst2_MC0_v1_1[1]), .ZN(Red_MCInst2_MC0_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC0_v0_1[1]), 
        .B(Red_MCInst2_MC0_v3_1[1]), .Z(Red_MCInst2_MC0_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC0_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC0_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[35]) );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC0_v2_1[2]), 
        .B(Red_MCInst2_MC0_v1_1[2]), .ZN(Red_MCInst2_MC0_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC0_v0_1[2]), 
        .B(Red_MCInst2_MC0_v3_1[2]), .Z(Red_MCInst2_MC0_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[21]) );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_2[0]), 
        .B(Red_MCInst2_MC0_v1_2[0]), .ZN(Red_MCInst2_MC0_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_2[0]), 
        .B(Red_MCInst2_MC0_v3_2[0]), .Z(Red_MCInst2_MC0_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC0_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC0_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[22]) );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC0_v2_2[1]), 
        .B(Red_MCInst2_MC0_v1_2[1]), .ZN(Red_MCInst2_MC0_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC0_v0_2[1]), 
        .B(Red_MCInst2_MC0_v3_2[1]), .Z(Red_MCInst2_MC0_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC0_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC0_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[23]) );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC0_v2_2[2]), 
        .B(Red_MCInst2_MC0_v1_2[2]), .ZN(Red_MCInst2_MC0_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), 
        .B(Red_MCInst2_MC0_v3_2[2]), .Z(Red_MCInst2_MC0_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[9]) );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC0_v2_3[0]), 
        .B(Red_MCInst2_MC0_v1_3[0]), .ZN(Red_MCInst2_MC0_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC0_v0_3[0]), 
        .B(Red_MCInst2_MC0_v3_3[0]), .Z(Red_MCInst2_MC0_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC0_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC0_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[10]) );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC0_v2_3[1]), 
        .B(Red_MCInst2_MC0_v1_3[1]), .ZN(Red_MCInst2_MC0_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC0_v0_3[1]), 
        .B(Red_MCInst2_MC0_v3_3[1]), .Z(Red_MCInst2_MC0_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC0_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC0_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[11]) );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC0_v2_3[2]), 
        .B(Red_MCInst2_MC0_v1_3[2]), .ZN(Red_MCInst2_MC0_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC0_v0_3[2]), 
        .B(Red_MCInst2_MC0_v3_3[2]), .Z(Red_MCInst2_MC0_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst2_MC1_U3 ( .A(ShiftRowsOutput2[24]), .Z(
        Red_MCInst2_MC1_v2_1[1]) );
  BUF_X1 Red_MCInst2_MC1_U2 ( .A(MCInst2_MC1_v1_3[2]), .Z(
        Red_MCInst2_MC1_v1_2[1]) );
  XOR2_X1 Red_MCInst2_MC1_v0_2Inst_0_U1 ( .A(MCInst2_MC1_v0_3[3]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(Red_MCInst2_MC1_v0_2[0]) );
  XOR2_X1 Red_MCInst2_MC1_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_2[2]), .Z(Red_MCInst2_MC1_v0_3[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC1_v1_0Inst_0_n3), 
        .B(MCInst2_MC1_v1_3[3]), .ZN(Red_MCInst2_MC1_v1_0[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_2[1]), .ZN(Red_MCInst2_MC1_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC1_v1_2Inst_0_U1 ( .A(Red_MCInst2_MC1_v1_2[1]), .B(
        Red_MCInst2_MC1_v1_1[2]), .Z(Red_MCInst2_MC1_v1_2[0]) );
  XOR2_X1 Red_MCInst2_MC1_v1_3Inst_0_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_2[1]), .Z(Red_MCInst2_MC1_v1_3[0]) );
  XOR2_X1 Red_MCInst2_MC1_v2_0Inst_0_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(Red_MCInst2_MC1_v2_0[0]) );
  XOR2_X1 Red_MCInst2_MC1_v2_1Inst_0_U1 ( .A(MCInst2_MC1_v2_0[2]), .B(
        MCInst2_MC1_v2_0[3]), .Z(Red_MCInst2_MC1_v2_1[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v2_2Inst_0_U2 ( .A(Red_MCInst2_MC1_v2_2Inst_0_n3), 
        .B(Red_MCInst2_MC1_v2_2[1]), .ZN(Red_MCInst2_MC1_v2_2[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v2_2Inst_0_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v2_0[2]), .ZN(Red_MCInst2_MC1_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v2_3Inst_0_U2 ( .A(Red_MCInst2_MC1_v2_3Inst_0_n3), 
        .B(Red_MCInst2_MC1_v2_2[1]), .ZN(Red_MCInst2_MC1_v2_3[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v2_3Inst_0_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v2_0[3]), .ZN(Red_MCInst2_MC1_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC1_v3_0Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_v3_0[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U3 ( .A(Red_MCInst2_MC1_v3_2Inst_0_n6), 
        .B(Red_MCInst2_MC1_v3_2Inst_0_n5), .ZN(Red_MCInst2_MC1_v3_2[0]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U2 ( .A(MCInst2_MC1_v3_0[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .ZN(Red_MCInst2_MC1_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC1_v3_3Inst_0_U1 ( .A(MCInst2_MC1_v3_0[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .Z(Red_MCInst2_MC1_v3_3[0]) );
  XOR2_X1 Red_MCInst2_MC1_v0_0Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), .B(
        Red_MCInst2_MC1_v0_1[0]), .Z(Red_MCInst2_MC1_v0_0[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v0_1Inst_1_U2 ( .A(Red_MCInst2_MC1_v0_1Inst_1_n3), 
        .B(Red_MCInst2_MC1_v0_1[0]), .ZN(Red_MCInst2_MC1_v0_1[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        MCInst2_MC1_v0_3[3]), .ZN(Red_MCInst2_MC1_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst2_MC1_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_2[2]), .Z(Red_MCInst2_MC1_v0_2[1]) );
  XOR2_X1 Red_MCInst2_MC1_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        MCInst2_MC1_v0_3[3]), .Z(Red_MCInst2_MC1_v0_3[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_1_U2 ( .A(Red_MCInst2_MC1_v1_0Inst_1_n3), 
        .B(Red_MCInst2_MC1_v1_1[2]), .ZN(Red_MCInst2_MC1_v1_0[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_2[1]), .ZN(Red_MCInst2_MC1_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v1_1Inst_1_U3 ( .A(Red_MCInst2_MC1_v1_1Inst_1_n6), 
        .B(Red_MCInst2_MC1_v1_1Inst_1_n5), .ZN(Red_MCInst2_MC1_v1_1[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_1Inst_1_U2 ( .A(MCInst2_MC1_v1_3[3]), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(Red_MCInst2_MC1_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC1_v1_1Inst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_2[1]), .Z(Red_MCInst2_MC1_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC1_v1_3Inst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        MCInst2_MC1_v1_3[3]), .Z(Red_MCInst2_MC1_v1_3[1]) );
  XOR2_X1 Red_MCInst2_MC1_v2_0Inst_1_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v2_0[3]), .Z(Red_MCInst2_MC1_v2_0[1]) );
  XOR2_X1 Red_MCInst2_MC1_v2_3Inst_1_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        Red_MCInst2_MC1_v2_2[1]), .Z(Red_MCInst2_MC1_v2_3[1]) );
  XOR2_X1 Red_MCInst2_MC1_v3_0Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[3]), .Z(Red_MCInst2_MC1_v3_0[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_1Inst_1_U3 ( .A(Red_MCInst2_MC1_v3_1Inst_1_n6), 
        .B(Red_MCInst2_MC1_v3_1Inst_1_n5), .ZN(Red_MCInst2_MC1_v3_1[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_1Inst_1_U2 ( .A(MCInst2_MC1_v3_0[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .ZN(Red_MCInst2_MC1_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC1_v3_1Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC1_v3_2Inst_1_U1 ( .A(Red_MCInst2_MC1_v3_3[2]), .B(
        MCInst2_MC1_v3_0[3]), .Z(Red_MCInst2_MC1_v3_2[1]) );
  XOR2_X1 Red_MCInst2_MC1_v3_3Inst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_v3_3[1]) );
  XNOR2_X1 Red_MCInst2_MC1_v0_0Inst_2_U2 ( .A(Red_MCInst2_MC1_v0_0Inst_2_n3), 
        .B(MCInst2_MC1_v0_3[3]), .ZN(Red_MCInst2_MC1_v0_0[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_2[2]), .ZN(Red_MCInst2_MC1_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst2_MC1_v0_1Inst_2_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_2[2]), .Z(Red_MCInst2_MC1_v0_1[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v0_3Inst_2_U3 ( .A(Red_MCInst2_MC1_v0_3Inst_2_n6), 
        .B(Red_MCInst2_MC1_v0_3Inst_2_n5), .ZN(Red_MCInst2_MC1_v0_3[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v0_3Inst_2_U2 ( .A(MCInst2_MC1_v0_3[3]), .B(
        Red_MCInst2_MC1_v0_1[0]), .ZN(Red_MCInst2_MC1_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC1_v0_3Inst_2_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), .B(
        Red_MCInst2_MC1_v0_2[2]), .Z(Red_MCInst2_MC1_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_2_U2 ( .A(Red_MCInst2_MC1_v1_0Inst_2_n3), 
        .B(Red_MCInst2_MC1_v1_1[2]), .ZN(Red_MCInst2_MC1_v1_0[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_2_U1 ( .A(Red_MCInst2_MC1_v1_2[1]), .B(
        MCInst2_MC1_v1_3[3]), .ZN(Red_MCInst2_MC1_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v1_2Inst_2_U2 ( .A(Red_MCInst2_MC1_v1_2Inst_2_n3), 
        .B(Red_MCInst2_MC1_v1_1[2]), .ZN(Red_MCInst2_MC1_v1_2[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_2Inst_2_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_2[1]), .ZN(Red_MCInst2_MC1_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC1_v1_3Inst_2_U3 ( .A(Red_MCInst2_MC1_v1_3Inst_2_n6), 
        .B(Red_MCInst2_MC1_v1_3Inst_2_n5), .ZN(Red_MCInst2_MC1_v1_3[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v1_3Inst_2_U2 ( .A(MCInst2_MC1_v1_3[3]), .B(
        Red_MCInst2_MC1_v1_1[2]), .ZN(Red_MCInst2_MC1_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC1_v1_3Inst_2_U1 ( .A(MCInst2_MC1_v1_0_0_), .B(
        Red_MCInst2_MC1_v1_2[1]), .Z(Red_MCInst2_MC1_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC1_v2_0Inst_2_U3 ( .A(Red_MCInst2_MC1_v2_0Inst_2_n6), 
        .B(Red_MCInst2_MC1_v2_0Inst_2_n5), .ZN(Red_MCInst2_MC1_v2_0[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v2_0Inst_2_U2 ( .A(MCInst2_MC1_v2_0[3]), .B(
        Red_MCInst2_MC1_v2_2[1]), .ZN(Red_MCInst2_MC1_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC1_v2_0Inst_2_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v2_0[2]), .Z(Red_MCInst2_MC1_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst2_MC1_v2_1Inst_2_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        Red_MCInst2_MC1_v2_2[1]), .Z(Red_MCInst2_MC1_v2_1[2]) );
  XOR2_X1 Red_MCInst2_MC1_v2_2Inst_2_U1 ( .A(MCInst2_MC1_v2_0[3]), .B(
        Red_MCInst2_MC1_v2_2[1]), .Z(Red_MCInst2_MC1_v2_2[2]) );
  XOR2_X1 Red_MCInst2_MC1_v2_3Inst_2_U1 ( .A(Red_MCInst2_MC1_v2_1[1]), .B(
        MCInst2_MC1_v2_0[3]), .Z(Red_MCInst2_MC1_v2_3[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_0Inst_2_U3 ( .A(Red_MCInst2_MC1_v3_0Inst_2_n6), 
        .B(Red_MCInst2_MC1_v3_0Inst_2_n5), .ZN(Red_MCInst2_MC1_v3_0[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_0Inst_2_U2 ( .A(MCInst2_MC1_v3_0[3]), .B(
        Red_MCInst2_MC1_v3_1[2]), .ZN(Red_MCInst2_MC1_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC1_v3_0Inst_2_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_2_U2 ( .A(Red_MCInst2_MC1_v3_2Inst_2_n3), 
        .B(Red_MCInst2_MC1_v3_1[2]), .ZN(Red_MCInst2_MC1_v3_2[2]) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_2_U1 ( .A(MCInst2_MC1_v3_2[3]), .B(
        MCInst2_MC1_v3_0[3]), .ZN(Red_MCInst2_MC1_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[42]) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_0[0]), 
        .B(Red_MCInst2_MC1_v1_0[0]), .ZN(Red_MCInst2_MC1_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), 
        .B(Red_MCInst2_MC1_v3_0[0]), .Z(Red_MCInst2_MC1_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC1_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC1_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[43]) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC1_v2_0[1]), 
        .B(Red_MCInst2_MC1_v1_0[1]), .ZN(Red_MCInst2_MC1_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC1_v0_0[1]), 
        .B(Red_MCInst2_MC1_v3_0[1]), .Z(Red_MCInst2_MC1_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC1_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC1_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[44]) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC1_v2_0[2]), 
        .B(Red_MCInst2_MC1_v1_0[2]), .ZN(Red_MCInst2_MC1_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC1_v0_0[2]), 
        .B(Red_MCInst2_MC1_v3_0[2]), .Z(Red_MCInst2_MC1_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[30]) );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_1[0]), 
        .B(Red_MCInst2_MC1_v1_2[1]), .ZN(Red_MCInst2_MC1_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_1[0]), 
        .B(Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC1_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC1_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[31]) );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC1_v2_1[1]), 
        .B(Red_MCInst2_MC1_v1_1[1]), .ZN(Red_MCInst2_MC1_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC1_v0_1[1]), 
        .B(Red_MCInst2_MC1_v3_1[1]), .Z(Red_MCInst2_MC1_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC1_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC1_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[32]) );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC1_v2_1[2]), 
        .B(Red_MCInst2_MC1_v1_1[2]), .ZN(Red_MCInst2_MC1_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC1_v0_1[2]), 
        .B(Red_MCInst2_MC1_v3_1[2]), .Z(Red_MCInst2_MC1_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[18]) );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_2[0]), 
        .B(Red_MCInst2_MC1_v1_2[0]), .ZN(Red_MCInst2_MC1_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_2[0]), 
        .B(Red_MCInst2_MC1_v3_2[0]), .Z(Red_MCInst2_MC1_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC1_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC1_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[19]) );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC1_v2_2[1]), 
        .B(Red_MCInst2_MC1_v1_2[1]), .ZN(Red_MCInst2_MC1_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC1_v0_2[1]), 
        .B(Red_MCInst2_MC1_v3_2[1]), .Z(Red_MCInst2_MC1_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC1_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC1_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[20]) );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC1_v2_2[2]), 
        .B(Red_MCInst2_MC1_v1_2[2]), .ZN(Red_MCInst2_MC1_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), 
        .B(Red_MCInst2_MC1_v3_2[2]), .Z(Red_MCInst2_MC1_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[6]) );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC1_v2_3[0]), 
        .B(Red_MCInst2_MC1_v1_3[0]), .ZN(Red_MCInst2_MC1_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC1_v0_3[0]), 
        .B(Red_MCInst2_MC1_v3_3[0]), .Z(Red_MCInst2_MC1_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC1_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC1_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[7]) );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC1_v2_3[1]), 
        .B(Red_MCInst2_MC1_v1_3[1]), .ZN(Red_MCInst2_MC1_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC1_v0_3[1]), 
        .B(Red_MCInst2_MC1_v3_3[1]), .Z(Red_MCInst2_MC1_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC1_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC1_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[8]) );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC1_v2_3[2]), 
        .B(Red_MCInst2_MC1_v1_3[2]), .ZN(Red_MCInst2_MC1_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC1_v0_3[2]), 
        .B(Red_MCInst2_MC1_v3_3[2]), .Z(Red_MCInst2_MC1_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst2_MC2_U3 ( .A(ShiftRowsOutput2[20]), .Z(
        Red_MCInst2_MC2_v2_1[1]) );
  BUF_X1 Red_MCInst2_MC2_U2 ( .A(MCInst2_MC2_v1_3[2]), .Z(
        Red_MCInst2_MC2_v1_2[1]) );
  XOR2_X1 Red_MCInst2_MC2_v0_2Inst_0_U1 ( .A(MCInst2_MC2_v0_3[3]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(Red_MCInst2_MC2_v0_2[0]) );
  XOR2_X1 Red_MCInst2_MC2_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_2[2]), .Z(Red_MCInst2_MC2_v0_3[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC2_v1_0Inst_0_n3), 
        .B(MCInst2_MC2_v1_3[3]), .ZN(Red_MCInst2_MC2_v1_0[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_2[1]), .ZN(Red_MCInst2_MC2_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC2_v1_2Inst_0_U1 ( .A(Red_MCInst2_MC2_v1_2[1]), .B(
        Red_MCInst2_MC2_v1_1[2]), .Z(Red_MCInst2_MC2_v1_2[0]) );
  XOR2_X1 Red_MCInst2_MC2_v1_3Inst_0_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_2[1]), .Z(Red_MCInst2_MC2_v1_3[0]) );
  XOR2_X1 Red_MCInst2_MC2_v2_0Inst_0_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(Red_MCInst2_MC2_v2_0[0]) );
  XOR2_X1 Red_MCInst2_MC2_v2_1Inst_0_U1 ( .A(MCInst2_MC2_v2_0[2]), .B(
        MCInst2_MC2_v2_0[3]), .Z(Red_MCInst2_MC2_v2_1[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v2_2Inst_0_U2 ( .A(Red_MCInst2_MC2_v2_2Inst_0_n3), 
        .B(Red_MCInst2_MC2_v2_2[1]), .ZN(Red_MCInst2_MC2_v2_2[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v2_2Inst_0_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v2_0[2]), .ZN(Red_MCInst2_MC2_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v2_3Inst_0_U2 ( .A(Red_MCInst2_MC2_v2_3Inst_0_n3), 
        .B(Red_MCInst2_MC2_v2_2[1]), .ZN(Red_MCInst2_MC2_v2_3[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v2_3Inst_0_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v2_0[3]), .ZN(Red_MCInst2_MC2_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC2_v3_0Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_v3_0[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U3 ( .A(Red_MCInst2_MC2_v3_2Inst_0_n6), 
        .B(Red_MCInst2_MC2_v3_2Inst_0_n5), .ZN(Red_MCInst2_MC2_v3_2[0]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U2 ( .A(MCInst2_MC2_v3_0[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .ZN(Red_MCInst2_MC2_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC2_v3_3Inst_0_U1 ( .A(MCInst2_MC2_v3_0[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .Z(Red_MCInst2_MC2_v3_3[0]) );
  XOR2_X1 Red_MCInst2_MC2_v0_0Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), .B(
        Red_MCInst2_MC2_v0_1[0]), .Z(Red_MCInst2_MC2_v0_0[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v0_1Inst_1_U2 ( .A(Red_MCInst2_MC2_v0_1Inst_1_n3), 
        .B(Red_MCInst2_MC2_v0_1[0]), .ZN(Red_MCInst2_MC2_v0_1[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        MCInst2_MC2_v0_3[3]), .ZN(Red_MCInst2_MC2_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst2_MC2_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_2[2]), .Z(Red_MCInst2_MC2_v0_2[1]) );
  XOR2_X1 Red_MCInst2_MC2_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        MCInst2_MC2_v0_3[3]), .Z(Red_MCInst2_MC2_v0_3[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_1_U2 ( .A(Red_MCInst2_MC2_v1_0Inst_1_n3), 
        .B(Red_MCInst2_MC2_v1_1[2]), .ZN(Red_MCInst2_MC2_v1_0[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_2[1]), .ZN(Red_MCInst2_MC2_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v1_1Inst_1_U3 ( .A(Red_MCInst2_MC2_v1_1Inst_1_n6), 
        .B(Red_MCInst2_MC2_v1_1Inst_1_n5), .ZN(Red_MCInst2_MC2_v1_1[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_1Inst_1_U2 ( .A(MCInst2_MC2_v1_3[3]), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(Red_MCInst2_MC2_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC2_v1_1Inst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_2[1]), .Z(Red_MCInst2_MC2_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC2_v1_3Inst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        MCInst2_MC2_v1_3[3]), .Z(Red_MCInst2_MC2_v1_3[1]) );
  XOR2_X1 Red_MCInst2_MC2_v2_0Inst_1_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v2_0[3]), .Z(Red_MCInst2_MC2_v2_0[1]) );
  XOR2_X1 Red_MCInst2_MC2_v2_3Inst_1_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        Red_MCInst2_MC2_v2_2[1]), .Z(Red_MCInst2_MC2_v2_3[1]) );
  XOR2_X1 Red_MCInst2_MC2_v3_0Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[3]), .Z(Red_MCInst2_MC2_v3_0[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_1Inst_1_U3 ( .A(Red_MCInst2_MC2_v3_1Inst_1_n6), 
        .B(Red_MCInst2_MC2_v3_1Inst_1_n5), .ZN(Red_MCInst2_MC2_v3_1[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_1Inst_1_U2 ( .A(MCInst2_MC2_v3_0[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .ZN(Red_MCInst2_MC2_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC2_v3_1Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC2_v3_2Inst_1_U1 ( .A(Red_MCInst2_MC2_v3_3[2]), .B(
        MCInst2_MC2_v3_0[3]), .Z(Red_MCInst2_MC2_v3_2[1]) );
  XOR2_X1 Red_MCInst2_MC2_v3_3Inst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_v3_3[1]) );
  XNOR2_X1 Red_MCInst2_MC2_v0_0Inst_2_U2 ( .A(Red_MCInst2_MC2_v0_0Inst_2_n3), 
        .B(MCInst2_MC2_v0_3[3]), .ZN(Red_MCInst2_MC2_v0_0[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_2[2]), .ZN(Red_MCInst2_MC2_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst2_MC2_v0_1Inst_2_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_2[2]), .Z(Red_MCInst2_MC2_v0_1[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v0_3Inst_2_U3 ( .A(Red_MCInst2_MC2_v0_3Inst_2_n6), 
        .B(Red_MCInst2_MC2_v0_3Inst_2_n5), .ZN(Red_MCInst2_MC2_v0_3[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v0_3Inst_2_U2 ( .A(MCInst2_MC2_v0_3[3]), .B(
        Red_MCInst2_MC2_v0_1[0]), .ZN(Red_MCInst2_MC2_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC2_v0_3Inst_2_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), .B(
        Red_MCInst2_MC2_v0_2[2]), .Z(Red_MCInst2_MC2_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_2_U2 ( .A(Red_MCInst2_MC2_v1_0Inst_2_n3), 
        .B(Red_MCInst2_MC2_v1_1[2]), .ZN(Red_MCInst2_MC2_v1_0[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_2_U1 ( .A(Red_MCInst2_MC2_v1_2[1]), .B(
        MCInst2_MC2_v1_3[3]), .ZN(Red_MCInst2_MC2_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v1_2Inst_2_U2 ( .A(Red_MCInst2_MC2_v1_2Inst_2_n3), 
        .B(Red_MCInst2_MC2_v1_1[2]), .ZN(Red_MCInst2_MC2_v1_2[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_2Inst_2_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_2[1]), .ZN(Red_MCInst2_MC2_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC2_v1_3Inst_2_U3 ( .A(Red_MCInst2_MC2_v1_3Inst_2_n6), 
        .B(Red_MCInst2_MC2_v1_3Inst_2_n5), .ZN(Red_MCInst2_MC2_v1_3[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v1_3Inst_2_U2 ( .A(MCInst2_MC2_v1_3[3]), .B(
        Red_MCInst2_MC2_v1_1[2]), .ZN(Red_MCInst2_MC2_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC2_v1_3Inst_2_U1 ( .A(MCInst2_MC2_v1_0_0_), .B(
        Red_MCInst2_MC2_v1_2[1]), .Z(Red_MCInst2_MC2_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC2_v2_0Inst_2_U3 ( .A(Red_MCInst2_MC2_v2_0Inst_2_n6), 
        .B(Red_MCInst2_MC2_v2_0Inst_2_n5), .ZN(Red_MCInst2_MC2_v2_0[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v2_0Inst_2_U2 ( .A(MCInst2_MC2_v2_0[3]), .B(
        Red_MCInst2_MC2_v2_2[1]), .ZN(Red_MCInst2_MC2_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC2_v2_0Inst_2_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v2_0[2]), .Z(Red_MCInst2_MC2_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst2_MC2_v2_1Inst_2_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        Red_MCInst2_MC2_v2_2[1]), .Z(Red_MCInst2_MC2_v2_1[2]) );
  XOR2_X1 Red_MCInst2_MC2_v2_2Inst_2_U1 ( .A(MCInst2_MC2_v2_0[3]), .B(
        Red_MCInst2_MC2_v2_2[1]), .Z(Red_MCInst2_MC2_v2_2[2]) );
  XOR2_X1 Red_MCInst2_MC2_v2_3Inst_2_U1 ( .A(Red_MCInst2_MC2_v2_1[1]), .B(
        MCInst2_MC2_v2_0[3]), .Z(Red_MCInst2_MC2_v2_3[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_0Inst_2_U3 ( .A(Red_MCInst2_MC2_v3_0Inst_2_n6), 
        .B(Red_MCInst2_MC2_v3_0Inst_2_n5), .ZN(Red_MCInst2_MC2_v3_0[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_0Inst_2_U2 ( .A(MCInst2_MC2_v3_0[3]), .B(
        Red_MCInst2_MC2_v3_1[2]), .ZN(Red_MCInst2_MC2_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC2_v3_0Inst_2_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_2_U2 ( .A(Red_MCInst2_MC2_v3_2Inst_2_n3), 
        .B(Red_MCInst2_MC2_v3_1[2]), .ZN(Red_MCInst2_MC2_v3_2[2]) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_2_U1 ( .A(MCInst2_MC2_v3_2[3]), .B(
        MCInst2_MC2_v3_0[3]), .ZN(Red_MCInst2_MC2_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[39]) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_0[0]), 
        .B(Red_MCInst2_MC2_v1_0[0]), .ZN(Red_MCInst2_MC2_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), 
        .B(Red_MCInst2_MC2_v3_0[0]), .Z(Red_MCInst2_MC2_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC2_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC2_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[40]) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC2_v2_0[1]), 
        .B(Red_MCInst2_MC2_v1_0[1]), .ZN(Red_MCInst2_MC2_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC2_v0_0[1]), 
        .B(Red_MCInst2_MC2_v3_0[1]), .Z(Red_MCInst2_MC2_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC2_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC2_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[41]) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC2_v2_0[2]), 
        .B(Red_MCInst2_MC2_v1_0[2]), .ZN(Red_MCInst2_MC2_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC2_v0_0[2]), 
        .B(Red_MCInst2_MC2_v3_0[2]), .Z(Red_MCInst2_MC2_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[27]) );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_1[0]), 
        .B(Red_MCInst2_MC2_v1_2[1]), .ZN(Red_MCInst2_MC2_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_1[0]), 
        .B(Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC2_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC2_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[28]) );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC2_v2_1[1]), 
        .B(Red_MCInst2_MC2_v1_1[1]), .ZN(Red_MCInst2_MC2_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC2_v0_1[1]), 
        .B(Red_MCInst2_MC2_v3_1[1]), .Z(Red_MCInst2_MC2_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC2_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC2_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[29]) );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC2_v2_1[2]), 
        .B(Red_MCInst2_MC2_v1_1[2]), .ZN(Red_MCInst2_MC2_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC2_v0_1[2]), 
        .B(Red_MCInst2_MC2_v3_1[2]), .Z(Red_MCInst2_MC2_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[15]) );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_2[0]), 
        .B(Red_MCInst2_MC2_v1_2[0]), .ZN(Red_MCInst2_MC2_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_2[0]), 
        .B(Red_MCInst2_MC2_v3_2[0]), .Z(Red_MCInst2_MC2_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC2_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC2_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[16]) );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC2_v2_2[1]), 
        .B(Red_MCInst2_MC2_v1_2[1]), .ZN(Red_MCInst2_MC2_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC2_v0_2[1]), 
        .B(Red_MCInst2_MC2_v3_2[1]), .Z(Red_MCInst2_MC2_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC2_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC2_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[17]) );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC2_v2_2[2]), 
        .B(Red_MCInst2_MC2_v1_2[2]), .ZN(Red_MCInst2_MC2_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), 
        .B(Red_MCInst2_MC2_v3_2[2]), .Z(Red_MCInst2_MC2_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[3]) );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC2_v2_3[0]), 
        .B(Red_MCInst2_MC2_v1_3[0]), .ZN(Red_MCInst2_MC2_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC2_v0_3[0]), 
        .B(Red_MCInst2_MC2_v3_3[0]), .Z(Red_MCInst2_MC2_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC2_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC2_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[4]) );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC2_v2_3[1]), 
        .B(Red_MCInst2_MC2_v1_3[1]), .ZN(Red_MCInst2_MC2_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC2_v0_3[1]), 
        .B(Red_MCInst2_MC2_v3_3[1]), .Z(Red_MCInst2_MC2_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC2_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC2_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[5]) );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC2_v2_3[2]), 
        .B(Red_MCInst2_MC2_v1_3[2]), .ZN(Red_MCInst2_MC2_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC2_v0_3[2]), 
        .B(Red_MCInst2_MC2_v3_3[2]), .Z(Red_MCInst2_MC2_r3Inst_XORInst_0_2_n8)
         );
  BUF_X1 Red_MCInst2_MC3_U3 ( .A(ShiftRowsOutput2[16]), .Z(
        Red_MCInst2_MC3_v2_1[1]) );
  BUF_X1 Red_MCInst2_MC3_U2 ( .A(MCInst2_MC3_v1_3[2]), .Z(
        Red_MCInst2_MC3_v1_2[1]) );
  XOR2_X1 Red_MCInst2_MC3_v0_2Inst_0_U1 ( .A(MCInst2_MC3_v0_3[3]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(Red_MCInst2_MC3_v0_2[0]) );
  XOR2_X1 Red_MCInst2_MC3_v0_3Inst_0_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_2[2]), .Z(Red_MCInst2_MC3_v0_3[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U2 ( .A(Red_MCInst2_MC3_v1_0Inst_0_n3), 
        .B(MCInst2_MC3_v1_3[3]), .ZN(Red_MCInst2_MC3_v1_0[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_2[1]), .ZN(Red_MCInst2_MC3_v1_0Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC3_v1_2Inst_0_U1 ( .A(Red_MCInst2_MC3_v1_2[1]), .B(
        Red_MCInst2_MC3_v1_1[2]), .Z(Red_MCInst2_MC3_v1_2[0]) );
  XOR2_X1 Red_MCInst2_MC3_v1_3Inst_0_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_2[1]), .Z(Red_MCInst2_MC3_v1_3[0]) );
  XOR2_X1 Red_MCInst2_MC3_v2_0Inst_0_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(Red_MCInst2_MC3_v2_0[0]) );
  XOR2_X1 Red_MCInst2_MC3_v2_1Inst_0_U1 ( .A(MCInst2_MC3_v2_0[2]), .B(
        MCInst2_MC3_v2_0[3]), .Z(Red_MCInst2_MC3_v2_1[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v2_2Inst_0_U2 ( .A(Red_MCInst2_MC3_v2_2Inst_0_n3), 
        .B(Red_MCInst2_MC3_v2_2[1]), .ZN(Red_MCInst2_MC3_v2_2[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v2_2Inst_0_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v2_0[2]), .ZN(Red_MCInst2_MC3_v2_2Inst_0_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v2_3Inst_0_U2 ( .A(Red_MCInst2_MC3_v2_3Inst_0_n3), 
        .B(Red_MCInst2_MC3_v2_2[1]), .ZN(Red_MCInst2_MC3_v2_3[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v2_3Inst_0_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v2_0[3]), .ZN(Red_MCInst2_MC3_v2_3Inst_0_n3) );
  XOR2_X1 Red_MCInst2_MC3_v3_0Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_v3_0[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U3 ( .A(Red_MCInst2_MC3_v3_2Inst_0_n6), 
        .B(Red_MCInst2_MC3_v3_2Inst_0_n5), .ZN(Red_MCInst2_MC3_v3_2[0]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U2 ( .A(MCInst2_MC3_v3_0[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .ZN(Red_MCInst2_MC3_v3_2Inst_0_n5) );
  XOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_v3_2Inst_0_n6) );
  XOR2_X1 Red_MCInst2_MC3_v3_3Inst_0_U1 ( .A(MCInst2_MC3_v3_0[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .Z(Red_MCInst2_MC3_v3_3[0]) );
  XOR2_X1 Red_MCInst2_MC3_v0_0Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), .B(
        Red_MCInst2_MC3_v0_1[0]), .Z(Red_MCInst2_MC3_v0_0[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v0_1Inst_1_U2 ( .A(Red_MCInst2_MC3_v0_1Inst_1_n3), 
        .B(Red_MCInst2_MC3_v0_1[0]), .ZN(Red_MCInst2_MC3_v0_1[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v0_1Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        MCInst2_MC3_v0_3[3]), .ZN(Red_MCInst2_MC3_v0_1Inst_1_n3) );
  XOR2_X1 Red_MCInst2_MC3_v0_2Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_2[2]), .Z(Red_MCInst2_MC3_v0_2[1]) );
  XOR2_X1 Red_MCInst2_MC3_v0_3Inst_1_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        MCInst2_MC3_v0_3[3]), .Z(Red_MCInst2_MC3_v0_3[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_1_U2 ( .A(Red_MCInst2_MC3_v1_0Inst_1_n3), 
        .B(Red_MCInst2_MC3_v1_1[2]), .ZN(Red_MCInst2_MC3_v1_0[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_2[1]), .ZN(Red_MCInst2_MC3_v1_0Inst_1_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v1_1Inst_1_U3 ( .A(Red_MCInst2_MC3_v1_1Inst_1_n6), 
        .B(Red_MCInst2_MC3_v1_1Inst_1_n5), .ZN(Red_MCInst2_MC3_v1_1[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_1Inst_1_U2 ( .A(MCInst2_MC3_v1_3[3]), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(Red_MCInst2_MC3_v1_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC3_v1_1Inst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_2[1]), .Z(Red_MCInst2_MC3_v1_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC3_v1_3Inst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        MCInst2_MC3_v1_3[3]), .Z(Red_MCInst2_MC3_v1_3[1]) );
  XOR2_X1 Red_MCInst2_MC3_v2_0Inst_1_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v2_0[3]), .Z(Red_MCInst2_MC3_v2_0[1]) );
  XOR2_X1 Red_MCInst2_MC3_v2_3Inst_1_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        Red_MCInst2_MC3_v2_2[1]), .Z(Red_MCInst2_MC3_v2_3[1]) );
  XOR2_X1 Red_MCInst2_MC3_v3_0Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[3]), .Z(Red_MCInst2_MC3_v3_0[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_1Inst_1_U3 ( .A(Red_MCInst2_MC3_v3_1Inst_1_n6), 
        .B(Red_MCInst2_MC3_v3_1Inst_1_n5), .ZN(Red_MCInst2_MC3_v3_1[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_1Inst_1_U2 ( .A(MCInst2_MC3_v3_0[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .ZN(Red_MCInst2_MC3_v3_1Inst_1_n5) );
  XOR2_X1 Red_MCInst2_MC3_v3_1Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_v3_1Inst_1_n6) );
  XOR2_X1 Red_MCInst2_MC3_v3_2Inst_1_U1 ( .A(Red_MCInst2_MC3_v3_3[2]), .B(
        MCInst2_MC3_v3_0[3]), .Z(Red_MCInst2_MC3_v3_2[1]) );
  XOR2_X1 Red_MCInst2_MC3_v3_3Inst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_v3_3[1]) );
  XNOR2_X1 Red_MCInst2_MC3_v0_0Inst_2_U2 ( .A(Red_MCInst2_MC3_v0_0Inst_2_n3), 
        .B(MCInst2_MC3_v0_3[3]), .ZN(Red_MCInst2_MC3_v0_0[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v0_0Inst_2_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_2[2]), .ZN(Red_MCInst2_MC3_v0_0Inst_2_n3) );
  XOR2_X1 Red_MCInst2_MC3_v0_1Inst_2_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_2[2]), .Z(Red_MCInst2_MC3_v0_1[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v0_3Inst_2_U3 ( .A(Red_MCInst2_MC3_v0_3Inst_2_n6), 
        .B(Red_MCInst2_MC3_v0_3Inst_2_n5), .ZN(Red_MCInst2_MC3_v0_3[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v0_3Inst_2_U2 ( .A(MCInst2_MC3_v0_3[3]), .B(
        Red_MCInst2_MC3_v0_1[0]), .ZN(Red_MCInst2_MC3_v0_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC3_v0_3Inst_2_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), .B(
        Red_MCInst2_MC3_v0_2[2]), .Z(Red_MCInst2_MC3_v0_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_2_U2 ( .A(Red_MCInst2_MC3_v1_0Inst_2_n3), 
        .B(Red_MCInst2_MC3_v1_1[2]), .ZN(Red_MCInst2_MC3_v1_0[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_2_U1 ( .A(Red_MCInst2_MC3_v1_2[1]), .B(
        MCInst2_MC3_v1_3[3]), .ZN(Red_MCInst2_MC3_v1_0Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v1_2Inst_2_U2 ( .A(Red_MCInst2_MC3_v1_2Inst_2_n3), 
        .B(Red_MCInst2_MC3_v1_1[2]), .ZN(Red_MCInst2_MC3_v1_2[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_2Inst_2_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_2[1]), .ZN(Red_MCInst2_MC3_v1_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC3_v1_3Inst_2_U3 ( .A(Red_MCInst2_MC3_v1_3Inst_2_n6), 
        .B(Red_MCInst2_MC3_v1_3Inst_2_n5), .ZN(Red_MCInst2_MC3_v1_3[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v1_3Inst_2_U2 ( .A(MCInst2_MC3_v1_3[3]), .B(
        Red_MCInst2_MC3_v1_1[2]), .ZN(Red_MCInst2_MC3_v1_3Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC3_v1_3Inst_2_U1 ( .A(MCInst2_MC3_v1_0_0_), .B(
        Red_MCInst2_MC3_v1_2[1]), .Z(Red_MCInst2_MC3_v1_3Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC3_v2_0Inst_2_U3 ( .A(Red_MCInst2_MC3_v2_0Inst_2_n6), 
        .B(Red_MCInst2_MC3_v2_0Inst_2_n5), .ZN(Red_MCInst2_MC3_v2_0[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v2_0Inst_2_U2 ( .A(MCInst2_MC3_v2_0[3]), .B(
        Red_MCInst2_MC3_v2_2[1]), .ZN(Red_MCInst2_MC3_v2_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC3_v2_0Inst_2_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v2_0[2]), .Z(Red_MCInst2_MC3_v2_0Inst_2_n6) );
  XOR2_X1 Red_MCInst2_MC3_v2_1Inst_2_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        Red_MCInst2_MC3_v2_2[1]), .Z(Red_MCInst2_MC3_v2_1[2]) );
  XOR2_X1 Red_MCInst2_MC3_v2_2Inst_2_U1 ( .A(MCInst2_MC3_v2_0[3]), .B(
        Red_MCInst2_MC3_v2_2[1]), .Z(Red_MCInst2_MC3_v2_2[2]) );
  XOR2_X1 Red_MCInst2_MC3_v2_3Inst_2_U1 ( .A(Red_MCInst2_MC3_v2_1[1]), .B(
        MCInst2_MC3_v2_0[3]), .Z(Red_MCInst2_MC3_v2_3[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_0Inst_2_U3 ( .A(Red_MCInst2_MC3_v3_0Inst_2_n6), 
        .B(Red_MCInst2_MC3_v3_0Inst_2_n5), .ZN(Red_MCInst2_MC3_v3_0[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_0Inst_2_U2 ( .A(MCInst2_MC3_v3_0[3]), .B(
        Red_MCInst2_MC3_v3_1[2]), .ZN(Red_MCInst2_MC3_v3_0Inst_2_n5) );
  XOR2_X1 Red_MCInst2_MC3_v3_0Inst_2_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_v3_0Inst_2_n6) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_2_U2 ( .A(Red_MCInst2_MC3_v3_2Inst_2_n3), 
        .B(Red_MCInst2_MC3_v3_1[2]), .ZN(Red_MCInst2_MC3_v3_2[2]) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_2_U1 ( .A(MCInst2_MC3_v3_2[3]), .B(
        MCInst2_MC3_v3_0[3]), .ZN(Red_MCInst2_MC3_v3_2Inst_2_n3) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[36]) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_0[0]), 
        .B(Red_MCInst2_MC3_v1_0[0]), .ZN(Red_MCInst2_MC3_r0Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), 
        .B(Red_MCInst2_MC3_v3_0[0]), .Z(Red_MCInst2_MC3_r0Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC3_r0Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC3_r0Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[37]) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC3_v2_0[1]), 
        .B(Red_MCInst2_MC3_v1_0[1]), .ZN(Red_MCInst2_MC3_r0Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC3_v0_0[1]), 
        .B(Red_MCInst2_MC3_v3_0[1]), .Z(Red_MCInst2_MC3_r0Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC3_r0Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC3_r0Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[38]) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC3_v2_0[2]), 
        .B(Red_MCInst2_MC3_v1_0[2]), .ZN(Red_MCInst2_MC3_r0Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC3_v0_0[2]), 
        .B(Red_MCInst2_MC3_v3_0[2]), .Z(Red_MCInst2_MC3_r0Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[24]) );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_1[0]), 
        .B(Red_MCInst2_MC3_v1_2[1]), .ZN(Red_MCInst2_MC3_r1Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_1[0]), 
        .B(Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_r1Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC3_r1Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC3_r1Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[25]) );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC3_v2_1[1]), 
        .B(Red_MCInst2_MC3_v1_1[1]), .ZN(Red_MCInst2_MC3_r1Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC3_v0_1[1]), 
        .B(Red_MCInst2_MC3_v3_1[1]), .Z(Red_MCInst2_MC3_r1Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC3_r1Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC3_r1Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[26]) );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC3_v2_1[2]), 
        .B(Red_MCInst2_MC3_v1_1[2]), .ZN(Red_MCInst2_MC3_r1Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC3_v0_1[2]), 
        .B(Red_MCInst2_MC3_v3_1[2]), .Z(Red_MCInst2_MC3_r1Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[12]) );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_2[0]), 
        .B(Red_MCInst2_MC3_v1_2[0]), .ZN(Red_MCInst2_MC3_r2Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_2[0]), 
        .B(Red_MCInst2_MC3_v3_2[0]), .Z(Red_MCInst2_MC3_r2Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC3_r2Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC3_r2Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[13]) );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC3_v2_2[1]), 
        .B(Red_MCInst2_MC3_v1_2[1]), .ZN(Red_MCInst2_MC3_r2Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC3_v0_2[1]), 
        .B(Red_MCInst2_MC3_v3_2[1]), .Z(Red_MCInst2_MC3_r2Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC3_r2Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC3_r2Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[14]) );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC3_v2_2[2]), 
        .B(Red_MCInst2_MC3_v1_2[2]), .ZN(Red_MCInst2_MC3_r2Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), 
        .B(Red_MCInst2_MC3_v3_2[2]), .Z(Red_MCInst2_MC3_r2Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U3 ( .A(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n8), .B(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n7), .ZN(Red_MC_output2[0]) );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U2 ( .A(Red_MCInst2_MC3_v2_3[0]), 
        .B(Red_MCInst2_MC3_v1_3[0]), .ZN(Red_MCInst2_MC3_r3Inst_XORInst_0_0_n7) );
  XOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U1 ( .A(Red_MCInst2_MC3_v0_3[0]), 
        .B(Red_MCInst2_MC3_v3_3[0]), .Z(Red_MCInst2_MC3_r3Inst_XORInst_0_0_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_1_U3 ( .A(
        Red_MCInst2_MC3_r3Inst_XORInst_0_1_n8), .B(
        Red_MCInst2_MC3_r3Inst_XORInst_0_1_n7), .ZN(Red_MC_output2[1]) );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_1_U2 ( .A(Red_MCInst2_MC3_v2_3[1]), 
        .B(Red_MCInst2_MC3_v1_3[1]), .ZN(Red_MCInst2_MC3_r3Inst_XORInst_0_1_n7) );
  XOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_1_U1 ( .A(Red_MCInst2_MC3_v0_3[1]), 
        .B(Red_MCInst2_MC3_v3_3[1]), .Z(Red_MCInst2_MC3_r3Inst_XORInst_0_1_n8)
         );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_2_U3 ( .A(
        Red_MCInst2_MC3_r3Inst_XORInst_0_2_n8), .B(
        Red_MCInst2_MC3_r3Inst_XORInst_0_2_n7), .ZN(Red_MC_output2[2]) );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_2_U2 ( .A(Red_MCInst2_MC3_v2_3[2]), 
        .B(Red_MCInst2_MC3_v1_3[2]), .ZN(Red_MCInst2_MC3_r3Inst_XORInst_0_2_n7) );
  XOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_2_U1 ( .A(Red_MCInst2_MC3_v0_3[2]), 
        .B(Red_MCInst2_MC3_v3_3[2]), .Z(Red_MCInst2_MC3_r3Inst_XORInst_0_2_n8)
         );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_0_LFInst_0_n3), .B(Key[2]), .ZN(Red_RoundKey[0]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_0_LFInst_1_n3), .B(Key[3]), .ZN(Red_RoundKey[1]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_1_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_0_LFInst_2_n3), .B(Key[3]), .ZN(Red_RoundKey[2]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_2_U1 ( .A(Key[1]), .B(Key[2]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_1_LFInst_0_n3), .B(Key[6]), .ZN(Red_RoundKey[3]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_1_LFInst_1_n3), .B(Key[7]), .ZN(Red_RoundKey[4]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_1_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_1_LFInst_2_n3), .B(Key[7]), .ZN(Red_RoundKey[5]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_2_U1 ( .A(Key[5]), .B(Key[6]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_2_LFInst_0_n3), .B(Key[10]), .ZN(Red_RoundKey[6])
         );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_2_LFInst_1_n3), .B(Key[11]), .ZN(Red_RoundKey[7])
         );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_1_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_2_LFInst_2_n3), .B(Key[11]), .ZN(Red_RoundKey[8])
         );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_2_U1 ( .A(Key[9]), .B(Key[10]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_3_LFInst_0_n3), .B(Key[14]), .ZN(Red_RoundKey[9])
         );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_3_LFInst_1_n3), .B(Key[15]), .ZN(Red_RoundKey[10])
         );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_1_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_3_LFInst_2_n3), .B(Key[15]), .ZN(Red_RoundKey[11])
         );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_2_U1 ( .A(Key[13]), .B(Key[14]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_4_LFInst_0_n3), .B(Key[18]), .ZN(Red_RoundKey[12])
         );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_4_LFInst_1_n3), .B(Key[19]), .ZN(Red_RoundKey[13])
         );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_1_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_4_LFInst_2_n3), .B(Key[19]), .ZN(Red_RoundKey[14])
         );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_2_U1 ( .A(Key[17]), .B(Key[18]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_5_LFInst_0_n3), .B(Key[22]), .ZN(Red_RoundKey[15])
         );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_5_LFInst_1_n3), .B(Key[23]), .ZN(Red_RoundKey[16])
         );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_1_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_5_LFInst_2_n3), .B(Key[23]), .ZN(Red_RoundKey[17])
         );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_2_U1 ( .A(Key[21]), .B(Key[22]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_6_LFInst_0_n3), .B(Key[26]), .ZN(Red_RoundKey[18])
         );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_6_LFInst_1_n3), .B(Key[27]), .ZN(Red_RoundKey[19])
         );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_1_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_6_LFInst_2_n3), .B(Key[27]), .ZN(Red_RoundKey[20])
         );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_2_U1 ( .A(Key[25]), .B(Key[26]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_7_LFInst_0_n3), .B(Key[30]), .ZN(Red_RoundKey[21])
         );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_7_LFInst_1_n3), .B(Key[31]), .ZN(Red_RoundKey[22])
         );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_1_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_7_LFInst_2_n3), .B(Key[31]), .ZN(Red_RoundKey[23])
         );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_2_U1 ( .A(Key[29]), .B(Key[30]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_8_LFInst_0_n3), .B(Key[34]), .ZN(Red_RoundKey[24])
         );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_8_LFInst_1_n3), .B(Key[35]), .ZN(Red_RoundKey[25])
         );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_1_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_8_LFInst_2_n3), .B(Key[35]), .ZN(Red_RoundKey[26])
         );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_2_U1 ( .A(Key[33]), .B(Key[34]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_9_LFInst_0_n3), .B(Key[38]), .ZN(Red_RoundKey[27])
         );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_9_LFInst_1_n3), .B(Key[39]), .ZN(Red_RoundKey[28])
         );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_1_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_9_LFInst_2_n3), .B(Key[39]), .ZN(Red_RoundKey[29])
         );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_2_U1 ( .A(Key[37]), .B(Key[38]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_10_LFInst_0_n3), .B(Key[42]), .ZN(Red_RoundKey[30])
         );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_10_LFInst_1_n3), .B(Key[43]), .ZN(Red_RoundKey[31])
         );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_1_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_10_LFInst_2_n3), .B(Key[43]), .ZN(Red_RoundKey[32])
         );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_2_U1 ( .A(Key[41]), .B(Key[42]), .ZN(
        Red_KeyInst_LFInst_10_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_11_LFInst_0_n3), .B(Key[46]), .ZN(Red_RoundKey[33])
         );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_11_LFInst_1_n3), .B(Key[47]), .ZN(Red_RoundKey[34])
         );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_1_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_11_LFInst_2_n3), .B(Key[47]), .ZN(Red_RoundKey[35])
         );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_2_U1 ( .A(Key[45]), .B(Key[46]), .ZN(
        Red_KeyInst_LFInst_11_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_12_LFInst_0_n3), .B(Key[50]), .ZN(Red_RoundKey[36])
         );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_12_LFInst_1_n3), .B(Key[51]), .ZN(Red_RoundKey[37])
         );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_1_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_12_LFInst_2_n3), .B(Key[51]), .ZN(Red_RoundKey[38])
         );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_2_U1 ( .A(Key[49]), .B(Key[50]), .ZN(
        Red_KeyInst_LFInst_12_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_13_LFInst_0_n3), .B(Key[54]), .ZN(Red_RoundKey[39])
         );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_13_LFInst_1_n3), .B(Key[55]), .ZN(Red_RoundKey[40])
         );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_1_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_13_LFInst_2_n3), .B(Key[55]), .ZN(Red_RoundKey[41])
         );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_2_U1 ( .A(Key[53]), .B(Key[54]), .ZN(
        Red_KeyInst_LFInst_13_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_14_LFInst_0_n3), .B(Key[58]), .ZN(Red_RoundKey[42])
         );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_14_LFInst_1_n3), .B(Key[59]), .ZN(Red_RoundKey[43])
         );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_1_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_14_LFInst_2_n3), .B(Key[59]), .ZN(Red_RoundKey[44])
         );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_2_U1 ( .A(Key[57]), .B(Key[58]), .ZN(
        Red_KeyInst_LFInst_14_LFInst_2_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_KeyInst_LFInst_15_LFInst_0_n3), .B(Key[62]), .ZN(Red_RoundKey[45])
         );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_0_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_KeyInst_LFInst_15_LFInst_1_n3), .B(Key[63]), .ZN(Red_RoundKey[46])
         );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_1_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_1_n3) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_KeyInst_LFInst_15_LFInst_2_n3), .B(Key[63]), .ZN(Red_RoundKey[47])
         );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_2_U1 ( .A(Key[61]), .B(Key[62]), .ZN(
        Red_KeyInst_LFInst_15_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_0_n3), .B(AddRoundKeyOutput[2]), .ZN(
        Red_SignaltoCheck[0]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_1_n3), .B(AddRoundKeyOutput[3]), .ZN(
        Red_SignaltoCheck[1]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_1_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_2_n3), .B(AddRoundKeyOutput[3]), .ZN(
        Red_SignaltoCheck[2]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[1]), 
        .B(AddRoundKeyOutput[2]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_0_n3), .B(AddRoundKeyOutput[6]), .ZN(
        Red_SignaltoCheck[3]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_1_n3), .B(AddRoundKeyOutput[7]), .ZN(
        Red_SignaltoCheck[4]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_1_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_2_n3), .B(AddRoundKeyOutput[7]), .ZN(
        Red_SignaltoCheck[5]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[5]), 
        .B(AddRoundKeyOutput[6]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_0_n3), .B(AddRoundKeyOutput[10]), .ZN(
        Red_SignaltoCheck[6]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_1_n3), .B(AddRoundKeyOutput[11]), .ZN(
        Red_SignaltoCheck[7]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_1_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_2_n3), .B(AddRoundKeyOutput[11]), .ZN(
        Red_SignaltoCheck[8]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_2_U1 ( .A(AddRoundKeyOutput[9]), 
        .B(AddRoundKeyOutput[10]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_0_n3), .B(AddRoundKeyOutput[14]), .ZN(
        Red_SignaltoCheck[9]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_1_n3), .B(AddRoundKeyOutput[15]), .ZN(
        Red_SignaltoCheck[10]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_1_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_2_n3), .B(AddRoundKeyOutput[15]), .ZN(
        Red_SignaltoCheck[11]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_2_U1 ( .A(AddRoundKeyOutput[13]), 
        .B(AddRoundKeyOutput[14]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_0_n3), .B(AddRoundKeyOutput[18]), .ZN(
        Red_SignaltoCheck[12]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_1_n3), .B(AddRoundKeyOutput[19]), .ZN(
        Red_SignaltoCheck[13]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_1_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_2_n3), .B(AddRoundKeyOutput[19]), .ZN(
        Red_SignaltoCheck[14]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_2_U1 ( .A(AddRoundKeyOutput[17]), 
        .B(AddRoundKeyOutput[18]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_0_n3), .B(AddRoundKeyOutput[22]), .ZN(
        Red_SignaltoCheck[15]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_1_n3), .B(AddRoundKeyOutput[23]), .ZN(
        Red_SignaltoCheck[16]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_1_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_2_n3), .B(AddRoundKeyOutput[23]), .ZN(
        Red_SignaltoCheck[17]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_2_U1 ( .A(AddRoundKeyOutput[21]), 
        .B(AddRoundKeyOutput[22]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_0_n3), .B(AddRoundKeyOutput[26]), .ZN(
        Red_SignaltoCheck[18]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_1_n3), .B(AddRoundKeyOutput[27]), .ZN(
        Red_SignaltoCheck[19]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_1_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_2_n3), .B(AddRoundKeyOutput[27]), .ZN(
        Red_SignaltoCheck[20]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_2_U1 ( .A(AddRoundKeyOutput[25]), 
        .B(AddRoundKeyOutput[26]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_0_n3), .B(AddRoundKeyOutput[30]), .ZN(
        Red_SignaltoCheck[21]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_1_n3), .B(AddRoundKeyOutput[31]), .ZN(
        Red_SignaltoCheck[22]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_1_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_2_n3), .B(AddRoundKeyOutput[31]), .ZN(
        Red_SignaltoCheck[23]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_2_U1 ( .A(AddRoundKeyOutput[29]), 
        .B(AddRoundKeyOutput[30]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_0_n3), .B(AddRoundKeyOutput[34]), .ZN(
        Red_SignaltoCheck[24]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_1_n3), .B(AddRoundKeyOutput[35]), .ZN(
        Red_SignaltoCheck[25]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_1_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_2_n3), .B(AddRoundKeyOutput[35]), .ZN(
        Red_SignaltoCheck[26]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_2_U1 ( .A(AddRoundKeyOutput[33]), 
        .B(AddRoundKeyOutput[34]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_0_n3), .B(AddRoundKeyOutput[38]), .ZN(
        Red_SignaltoCheck[27]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_1_n3), .B(AddRoundKeyOutput[39]), .ZN(
        Red_SignaltoCheck[28]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_1_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_2_n3), .B(AddRoundKeyOutput[39]), .ZN(
        Red_SignaltoCheck[29]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_2_U1 ( .A(AddRoundKeyOutput[37]), 
        .B(AddRoundKeyOutput[38]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_0_n3), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_1_n3), .B(AddRoundKeyOutput[43]), 
        .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_1_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_2_n3), .B(AddRoundKeyOutput[43]), 
        .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_2_U1 ( .A(AddRoundKeyOutput[41]), 
        .B(AddRoundKeyOutput[42]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_0_n3), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_1_n3), .B(AddRoundKeyOutput[47]), 
        .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_1_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_2_n3), .B(AddRoundKeyOutput[47]), 
        .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[45]), 
        .B(AddRoundKeyOutput[46]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_0_n3), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_1_n3), .B(AddRoundKeyOutput[51]), 
        .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_1_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_2_n3), .B(AddRoundKeyOutput[51]), 
        .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_2_U1 ( .A(AddRoundKeyOutput[49]), 
        .B(AddRoundKeyOutput[50]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_0_n3), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_1_n3), .B(AddRoundKeyOutput[55]), 
        .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_1_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_2_n3), .B(AddRoundKeyOutput[55]), 
        .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[53]), 
        .B(AddRoundKeyOutput[54]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_0_n3), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_1_n3), .B(AddRoundKeyOutput[59]), 
        .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_1_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_2_n3), .B(AddRoundKeyOutput[59]), 
        .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_2_U1 ( .A(AddRoundKeyOutput[57]), 
        .B(AddRoundKeyOutput[58]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_0_n3), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_1_n3), .B(AddRoundKeyOutput[63]), 
        .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_1_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_2_n3), .B(AddRoundKeyOutput[63]), 
        .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_2_U1 ( .A(AddRoundKeyOutput[61]), 
        .B(AddRoundKeyOutput[62]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_2_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_0_n3), .B(Ciphertext[2]), .ZN(
        Red_SignaltoCheck[48]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U1 ( .A(Ciphertext[0]), .B(
        Ciphertext[1]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_1_n3), .B(Ciphertext[3]), .ZN(
        Red_SignaltoCheck[49]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_1_U1 ( .A(Ciphertext[0]), .B(
        Ciphertext[1]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_2_n3), .B(Ciphertext[3]), .ZN(
        Red_SignaltoCheck[50]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_2_U1 ( .A(Ciphertext[1]), .B(
        Ciphertext[2]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_0_n3), .B(Ciphertext[6]), .ZN(
        Red_SignaltoCheck[51]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U1 ( .A(Ciphertext[4]), .B(
        Ciphertext[5]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_1_n3), .B(Ciphertext[7]), .ZN(
        Red_SignaltoCheck[52]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_1_U1 ( .A(Ciphertext[4]), .B(
        Ciphertext[5]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_2_n3), .B(Ciphertext[7]), .ZN(
        Red_SignaltoCheck[53]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_2_U1 ( .A(Ciphertext[5]), .B(
        Ciphertext[6]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_0_n3), .B(Ciphertext[10]), .ZN(
        Red_SignaltoCheck[54]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U1 ( .A(Ciphertext[8]), .B(
        Ciphertext[9]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_1_n3), .B(Ciphertext[11]), .ZN(
        Red_SignaltoCheck[55]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_1_U1 ( .A(Ciphertext[8]), .B(
        Ciphertext[9]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_2_n3), .B(Ciphertext[11]), .ZN(
        Red_SignaltoCheck[56]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_2_U1 ( .A(Ciphertext[9]), .B(
        Ciphertext[10]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_0_n3), .B(Ciphertext[14]), .ZN(
        Red_SignaltoCheck[57]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U1 ( .A(Ciphertext[12]), .B(
        Ciphertext[13]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_1_n3), .B(Ciphertext[15]), .ZN(
        Red_SignaltoCheck[58]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_1_U1 ( .A(Ciphertext[12]), .B(
        Ciphertext[13]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_2_n3), .B(Ciphertext[15]), .ZN(
        Red_SignaltoCheck[59]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_2_U1 ( .A(Ciphertext[13]), .B(
        Ciphertext[14]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_0_n3), .B(Ciphertext[18]), .ZN(
        Red_SignaltoCheck[60]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U1 ( .A(Ciphertext[16]), .B(
        Ciphertext[17]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_1_n3), .B(Ciphertext[19]), .ZN(
        Red_SignaltoCheck[61]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_1_U1 ( .A(Ciphertext[16]), .B(
        Ciphertext[17]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_2_n3), .B(Ciphertext[19]), .ZN(
        Red_SignaltoCheck[62]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_2_U1 ( .A(Ciphertext[17]), .B(
        Ciphertext[18]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_0_n3), .B(Ciphertext[22]), .ZN(
        Red_SignaltoCheck[63]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U1 ( .A(Ciphertext[20]), .B(
        Ciphertext[21]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_1_n3), .B(Ciphertext[23]), .ZN(
        Red_SignaltoCheck[64]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_1_U1 ( .A(Ciphertext[20]), .B(
        Ciphertext[21]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_2_n3), .B(Ciphertext[23]), .ZN(
        Red_SignaltoCheck[65]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_2_U1 ( .A(Ciphertext[21]), .B(
        Ciphertext[22]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_0_n3), .B(Ciphertext[26]), .ZN(
        Red_SignaltoCheck[66]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U1 ( .A(Ciphertext[24]), .B(
        Ciphertext[25]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_1_n3), .B(Ciphertext[27]), .ZN(
        Red_SignaltoCheck[67]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_1_U1 ( .A(Ciphertext[24]), .B(
        Ciphertext[25]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_2_n3), .B(Ciphertext[27]), .ZN(
        Red_SignaltoCheck[68]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_2_U1 ( .A(Ciphertext[25]), .B(
        Ciphertext[26]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_0_n3), .B(Ciphertext[30]), .ZN(
        Red_SignaltoCheck[69]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U1 ( .A(Ciphertext[28]), .B(
        Ciphertext[29]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_1_n3), .B(Ciphertext[31]), .ZN(
        Red_SignaltoCheck[70]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_1_U1 ( .A(Ciphertext[28]), .B(
        Ciphertext[29]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_2_n3), .B(Ciphertext[31]), .ZN(
        Red_SignaltoCheck[71]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_2_U1 ( .A(Ciphertext[29]), .B(
        Ciphertext[30]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_0_n3), .B(Ciphertext[34]), .ZN(
        Red_SignaltoCheck[72]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U1 ( .A(Ciphertext[32]), .B(
        Ciphertext[33]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_1_n3), .B(Ciphertext[35]), .ZN(
        Red_SignaltoCheck[73]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_1_U1 ( .A(Ciphertext[32]), .B(
        Ciphertext[33]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_2_n3), .B(Ciphertext[35]), .ZN(
        Red_SignaltoCheck[74]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_2_U1 ( .A(Ciphertext[33]), .B(
        Ciphertext[34]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_0_n3), .B(Ciphertext[38]), .ZN(
        Red_SignaltoCheck[75]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U1 ( .A(Ciphertext[36]), .B(
        Ciphertext[37]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_1_n3), .B(Ciphertext[39]), .ZN(
        Red_SignaltoCheck[76]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_1_U1 ( .A(Ciphertext[36]), .B(
        Ciphertext[37]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_2_n3), .B(Ciphertext[39]), .ZN(
        Red_SignaltoCheck[77]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_2_U1 ( .A(Ciphertext[37]), .B(
        Ciphertext[38]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_0_n3), .B(Ciphertext[42]), .ZN(
        Red_SignaltoCheck[78]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U1 ( .A(Ciphertext[40]), .B(
        Ciphertext[41]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_1_n3), .B(Ciphertext[43]), .ZN(
        Red_SignaltoCheck[79]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_1_U1 ( .A(Ciphertext[40]), .B(
        Ciphertext[41]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_2_n3), .B(Ciphertext[43]), .ZN(
        Red_SignaltoCheck[80]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_2_U1 ( .A(Ciphertext[41]), .B(
        Ciphertext[42]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_0_n3), .B(Ciphertext[46]), .ZN(
        Red_SignaltoCheck[81]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U1 ( .A(Ciphertext[44]), .B(
        Ciphertext[45]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_1_n3), .B(Ciphertext[47]), .ZN(
        Red_SignaltoCheck[82]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_1_U1 ( .A(Ciphertext[44]), .B(
        Ciphertext[45]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_2_n3), .B(Ciphertext[47]), .ZN(
        Red_SignaltoCheck[83]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_2_U1 ( .A(Ciphertext[45]), .B(
        Ciphertext[46]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_0_n3), .B(Ciphertext[50]), .ZN(
        Red_SignaltoCheck[84]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U1 ( .A(Ciphertext[48]), .B(
        Ciphertext[49]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_1_n3), .B(Ciphertext[51]), .ZN(
        Red_SignaltoCheck[85]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_1_U1 ( .A(Ciphertext[48]), .B(
        Ciphertext[49]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_2_n3), .B(Ciphertext[51]), .ZN(
        Red_SignaltoCheck[86]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_2_U1 ( .A(Ciphertext[49]), .B(
        Ciphertext[50]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_0_n3), .B(Ciphertext[54]), .ZN(
        Red_SignaltoCheck[87]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U1 ( .A(Ciphertext[52]), .B(
        Ciphertext[53]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_1_n3), .B(Ciphertext[55]), .ZN(
        Red_SignaltoCheck[88]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_1_U1 ( .A(Ciphertext[52]), .B(
        Ciphertext[53]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_2_n3), .B(Ciphertext[55]), .ZN(
        Red_SignaltoCheck[89]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_2_U1 ( .A(Ciphertext[53]), .B(
        Ciphertext[54]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_0_n3), .B(Ciphertext[58]), .ZN(
        Red_SignaltoCheck[90]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U1 ( .A(Ciphertext[56]), .B(
        Ciphertext[57]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_1_n3), .B(Ciphertext[59]), .ZN(
        Red_SignaltoCheck[91]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_1_U1 ( .A(Ciphertext[56]), .B(
        Ciphertext[57]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_2_n3), .B(Ciphertext[59]), .ZN(
        Red_SignaltoCheck[92]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_2_U1 ( .A(Ciphertext[57]), .B(
        Ciphertext[58]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_0_n3), .B(Ciphertext[62]), .ZN(
        Red_SignaltoCheck[93]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U1 ( .A(Ciphertext[60]), .B(
        Ciphertext[61]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_1_n3), .B(Ciphertext[63]), .ZN(
        Red_SignaltoCheck[94]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_1_U1 ( .A(Ciphertext[60]), .B(
        Ciphertext[61]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_2_n3), .B(Ciphertext[63]), .ZN(
        Red_SignaltoCheck[95]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_2_U1 ( .A(Ciphertext[61]), .B(
        Ciphertext[62]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_0_n3), .B(MCInst2_MC3_v3_0[3]), .ZN(
        Red_SignaltoCheck[96]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U1 ( .A(MCInst2_MC3_v3_2[3]), 
        .B(Red_MCInst2_MC3_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_1_n3), .B(Red_MCInst2_MC3_v3_1[2]), 
        .ZN(Red_SignaltoCheck[97]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_1_U1 ( .A(MCInst2_MC3_v3_2[3]), 
        .B(Red_MCInst2_MC3_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_2_n3), .B(Red_MCInst2_MC3_v3_1[2]), 
        .ZN(Red_SignaltoCheck[98]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_2_U1 ( .A(Red_MCInst2_MC3_v3_3[2]), 
        .B(MCInst2_MC3_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_0_n3), .B(MCInst2_MC2_v3_0[3]), .ZN(
        Red_SignaltoCheck[99]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U1 ( .A(MCInst2_MC2_v3_2[3]), 
        .B(Red_MCInst2_MC2_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_1_n3), .B(Red_MCInst2_MC2_v3_1[2]), 
        .ZN(Red_SignaltoCheck[100]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_1_U1 ( .A(MCInst2_MC2_v3_2[3]), 
        .B(Red_MCInst2_MC2_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_2_n3), .B(Red_MCInst2_MC2_v3_1[2]), 
        .ZN(Red_SignaltoCheck[101]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_2_U1 ( .A(Red_MCInst2_MC2_v3_3[2]), 
        .B(MCInst2_MC2_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_0_n3), .B(MCInst2_MC1_v3_0[3]), .ZN(
        Red_SignaltoCheck[102]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U1 ( .A(MCInst2_MC1_v3_2[3]), 
        .B(Red_MCInst2_MC1_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_1_n3), .B(Red_MCInst2_MC1_v3_1[2]), 
        .ZN(Red_SignaltoCheck[103]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_1_U1 ( .A(MCInst2_MC1_v3_2[3]), 
        .B(Red_MCInst2_MC1_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_2_n3), .B(Red_MCInst2_MC1_v3_1[2]), 
        .ZN(Red_SignaltoCheck[104]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_2_U1 ( .A(Red_MCInst2_MC1_v3_3[2]), 
        .B(MCInst2_MC1_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_0_n3), .B(MCInst2_MC0_v3_0[3]), .ZN(
        Red_SignaltoCheck[105]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U1 ( .A(MCInst2_MC0_v3_2[3]), 
        .B(Red_MCInst2_MC0_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_1_n3), .B(Red_MCInst2_MC0_v3_1[2]), 
        .ZN(Red_SignaltoCheck[106]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_1_U1 ( .A(MCInst2_MC0_v3_2[3]), 
        .B(Red_MCInst2_MC0_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_2_n3), .B(Red_MCInst2_MC0_v3_1[2]), 
        .ZN(Red_SignaltoCheck[107]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_2_U1 ( .A(Red_MCInst2_MC0_v3_3[2]), 
        .B(MCInst2_MC0_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_0_n3), .B(MCInst2_MC3_v2_0[3]), .ZN(
        Red_SignaltoCheck[108]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U1 ( .A(ShiftRowsOutput2[16]), 
        .B(MCInst2_MC3_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_1_n3), .B(Red_MCInst2_MC3_v2_2[1]), 
        .ZN(Red_SignaltoCheck[109]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_1_U1 ( .A(ShiftRowsOutput2[16]), 
        .B(MCInst2_MC3_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_2_n3), .B(Red_MCInst2_MC3_v2_2[1]), 
        .ZN(Red_SignaltoCheck[110]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_2_U1 ( .A(MCInst2_MC3_v2_0[2]), 
        .B(MCInst2_MC3_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_0_n3), .B(MCInst2_MC2_v2_0[3]), .ZN(
        Red_SignaltoCheck[111]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U1 ( .A(ShiftRowsOutput2[20]), 
        .B(MCInst2_MC2_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_1_n3), .B(Red_MCInst2_MC2_v2_2[1]), 
        .ZN(Red_SignaltoCheck[112]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_1_U1 ( .A(ShiftRowsOutput2[20]), 
        .B(MCInst2_MC2_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_2_n3), .B(Red_MCInst2_MC2_v2_2[1]), 
        .ZN(Red_SignaltoCheck[113]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_2_U1 ( .A(MCInst2_MC2_v2_0[2]), 
        .B(MCInst2_MC2_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_0_n3), .B(MCInst2_MC1_v2_0[3]), .ZN(
        Red_SignaltoCheck[114]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U1 ( .A(ShiftRowsOutput2[24]), 
        .B(MCInst2_MC1_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_1_n3), .B(Red_MCInst2_MC1_v2_2[1]), 
        .ZN(Red_SignaltoCheck[115]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_1_U1 ( .A(ShiftRowsOutput2[24]), 
        .B(MCInst2_MC1_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_2_n3), .B(Red_MCInst2_MC1_v2_2[1]), 
        .ZN(Red_SignaltoCheck[116]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_2_U1 ( .A(MCInst2_MC1_v2_0[2]), 
        .B(MCInst2_MC1_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_0_n3), .B(MCInst2_MC0_v2_0[3]), .ZN(
        Red_SignaltoCheck[117]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U1 ( .A(ShiftRowsOutput2[28]), 
        .B(MCInst2_MC0_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_1_n3), .B(Red_MCInst2_MC0_v2_2[1]), 
        .ZN(Red_SignaltoCheck[118]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_1_U1 ( .A(ShiftRowsOutput2[28]), 
        .B(MCInst2_MC0_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_2_n3), .B(Red_MCInst2_MC0_v2_2[1]), 
        .ZN(Red_SignaltoCheck[119]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_2_U1 ( .A(MCInst2_MC0_v2_0[2]), 
        .B(MCInst2_MC0_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_0_n3), .B(MCInst2_MC3_v1_3[3]), .ZN(
        Red_SignaltoCheck[120]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U1 ( .A(MCInst2_MC3_v1_0_0_), 
        .B(MCInst2_MC3_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_1_n3), .B(Red_MCInst2_MC3_v1_1[2]), 
        .ZN(Red_SignaltoCheck[121]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_1_U1 ( .A(MCInst2_MC3_v1_0_0_), 
        .B(MCInst2_MC3_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_2_n3), .B(Red_MCInst2_MC3_v1_1[2]), 
        .ZN(Red_SignaltoCheck[122]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_2_U1 ( .A(MCInst2_MC3_v1_3[2]), 
        .B(MCInst2_MC3_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_0_n3), .B(MCInst2_MC2_v1_3[3]), .ZN(
        Red_SignaltoCheck[123]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U1 ( .A(MCInst2_MC2_v1_0_0_), 
        .B(MCInst2_MC2_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_1_n3), .B(Red_MCInst2_MC2_v1_1[2]), 
        .ZN(Red_SignaltoCheck[124]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_1_U1 ( .A(MCInst2_MC2_v1_0_0_), 
        .B(MCInst2_MC2_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_2_n3), .B(Red_MCInst2_MC2_v1_1[2]), 
        .ZN(Red_SignaltoCheck[125]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_2_U1 ( .A(MCInst2_MC2_v1_3[2]), 
        .B(MCInst2_MC2_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_0_n3), .B(MCInst2_MC1_v1_3[3]), .ZN(
        Red_SignaltoCheck[126]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U1 ( .A(MCInst2_MC1_v1_0_0_), 
        .B(MCInst2_MC1_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_1_n3), .B(Red_MCInst2_MC1_v1_1[2]), 
        .ZN(Red_SignaltoCheck[127]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_1_U1 ( .A(MCInst2_MC1_v1_0_0_), 
        .B(MCInst2_MC1_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_2_n3), .B(Red_MCInst2_MC1_v1_1[2]), 
        .ZN(Red_SignaltoCheck[128]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_2_U1 ( .A(MCInst2_MC1_v1_3[2]), 
        .B(MCInst2_MC1_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_0_n3), .B(MCInst2_MC0_v1_3[3]), .ZN(
        Red_SignaltoCheck[129]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U1 ( .A(MCInst2_MC0_v1_0_0_), 
        .B(MCInst2_MC0_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_1_n3), .B(Red_MCInst2_MC0_v1_1[2]), 
        .ZN(Red_SignaltoCheck[130]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_1_U1 ( .A(MCInst2_MC0_v1_0_0_), 
        .B(MCInst2_MC0_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_2_n3), .B(Red_MCInst2_MC0_v1_1[2]), 
        .ZN(Red_SignaltoCheck[131]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_2_U1 ( .A(MCInst2_MC0_v1_3[2]), 
        .B(MCInst2_MC0_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_0_n3), .B(MCInst2_MC3_v0_3[3]), .ZN(
        Red_SignaltoCheck[132]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), 
        .B(Red_MCInst2_MC3_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_1_n3), .B(Red_MCInst2_MC3_v0_1[0]), 
        .ZN(Red_SignaltoCheck[133]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_1_U1 ( .A(Red_MCInst2_MC3_v0_0[0]), 
        .B(Red_MCInst2_MC3_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_2_n3), .B(Red_MCInst2_MC3_v0_1[0]), 
        .ZN(Red_SignaltoCheck[134]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_2_U1 ( .A(Red_MCInst2_MC3_v0_2[2]), 
        .B(MCInst2_MC3_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_0_n3), .B(MCInst2_MC2_v0_3[3]), .ZN(
        Red_SignaltoCheck[135]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), 
        .B(Red_MCInst2_MC2_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_1_n3), .B(Red_MCInst2_MC2_v0_1[0]), 
        .ZN(Red_SignaltoCheck[136]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_1_U1 ( .A(Red_MCInst2_MC2_v0_0[0]), 
        .B(Red_MCInst2_MC2_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_2_n3), .B(Red_MCInst2_MC2_v0_1[0]), 
        .ZN(Red_SignaltoCheck[137]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_2_U1 ( .A(Red_MCInst2_MC2_v0_2[2]), 
        .B(MCInst2_MC2_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_0_n3), .B(MCInst2_MC1_v0_3[3]), .ZN(
        Red_SignaltoCheck[138]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), 
        .B(Red_MCInst2_MC1_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_1_n3), .B(Red_MCInst2_MC1_v0_1[0]), 
        .ZN(Red_SignaltoCheck[139]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_1_U1 ( .A(Red_MCInst2_MC1_v0_0[0]), 
        .B(Red_MCInst2_MC1_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_2_n3), .B(Red_MCInst2_MC1_v0_1[0]), 
        .ZN(Red_SignaltoCheck[140]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_2_U1 ( .A(Red_MCInst2_MC1_v0_2[2]), 
        .B(MCInst2_MC1_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_0_n3), .B(MCInst2_MC0_v0_3[3]), .ZN(
        Red_SignaltoCheck[141]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), 
        .B(Red_MCInst2_MC0_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_1_n3), .B(Red_MCInst2_MC0_v0_1[0]), 
        .ZN(Red_SignaltoCheck[142]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_1_U1 ( .A(Red_MCInst2_MC0_v0_0[0]), 
        .B(Red_MCInst2_MC0_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_2_n3), .B(Red_MCInst2_MC0_v0_1[0]), 
        .ZN(Red_SignaltoCheck[143]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_2_U1 ( .A(Red_MCInst2_MC0_v0_2[2]), 
        .B(MCInst2_MC0_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_48_LFInst_0_n3), .B(SubCellInput2[2]), .ZN(
        Red_SignaltoCheck[144]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U1 ( .A(SubCellInput2[0]), .B(
        SubCellInput2[1]), .ZN(Red_ToCheckInst_LFInst_48_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_48_LFInst_1_n3), .B(SubCellInput2[3]), .ZN(
        Red_SignaltoCheck[145]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_1_U1 ( .A(SubCellInput2[0]), .B(
        SubCellInput2[1]), .ZN(Red_ToCheckInst_LFInst_48_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_48_LFInst_2_n3), .B(SubCellInput2[3]), .ZN(
        Red_SignaltoCheck[146]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_2_U1 ( .A(SubCellInput2[1]), .B(
        SubCellInput2[2]), .ZN(Red_ToCheckInst_LFInst_48_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_49_LFInst_0_n3), .B(SubCellInput2[6]), .ZN(
        Red_SignaltoCheck[147]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U1 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[5]), .ZN(Red_ToCheckInst_LFInst_49_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_49_LFInst_1_n3), .B(SubCellInput2[7]), .ZN(
        Red_SignaltoCheck[148]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_1_U1 ( .A(SubCellInput2[4]), .B(
        SubCellInput2[5]), .ZN(Red_ToCheckInst_LFInst_49_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_49_LFInst_2_n3), .B(SubCellInput2[7]), .ZN(
        Red_SignaltoCheck[149]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_2_U1 ( .A(SubCellInput2[5]), .B(
        SubCellInput2[6]), .ZN(Red_ToCheckInst_LFInst_49_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_50_LFInst_0_n3), .B(SubCellInput2[10]), .ZN(
        Red_SignaltoCheck[150]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U1 ( .A(SubCellInput2[8]), .B(
        SubCellInput2[9]), .ZN(Red_ToCheckInst_LFInst_50_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_50_LFInst_1_n3), .B(SubCellInput2[11]), .ZN(
        Red_SignaltoCheck[151]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_1_U1 ( .A(SubCellInput2[8]), .B(
        SubCellInput2[9]), .ZN(Red_ToCheckInst_LFInst_50_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_50_LFInst_2_n3), .B(SubCellInput2[11]), .ZN(
        Red_SignaltoCheck[152]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_2_U1 ( .A(SubCellInput2[9]), .B(
        SubCellInput2[10]), .ZN(Red_ToCheckInst_LFInst_50_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_51_LFInst_0_n3), .B(SubCellInput2[14]), .ZN(
        Red_SignaltoCheck[153]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U1 ( .A(SubCellInput2[12]), .B(
        SubCellInput2[13]), .ZN(Red_ToCheckInst_LFInst_51_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_51_LFInst_1_n3), .B(SubCellInput2[15]), .ZN(
        Red_SignaltoCheck[154]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_1_U1 ( .A(SubCellInput2[12]), .B(
        SubCellInput2[13]), .ZN(Red_ToCheckInst_LFInst_51_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_51_LFInst_2_n3), .B(SubCellInput2[15]), .ZN(
        Red_SignaltoCheck[155]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_2_U1 ( .A(SubCellInput2[13]), .B(
        SubCellInput2[14]), .ZN(Red_ToCheckInst_LFInst_51_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_52_LFInst_0_n3), .B(SubCellInput2[18]), .ZN(
        Red_SignaltoCheck[156]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U1 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[17]), .ZN(Red_ToCheckInst_LFInst_52_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_52_LFInst_1_n3), .B(SubCellInput2[19]), .ZN(
        Red_SignaltoCheck[157]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_1_U1 ( .A(SubCellInput2[16]), .B(
        SubCellInput2[17]), .ZN(Red_ToCheckInst_LFInst_52_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_52_LFInst_2_n3), .B(SubCellInput2[19]), .ZN(
        Red_SignaltoCheck[158]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_2_U1 ( .A(SubCellInput2[17]), .B(
        SubCellInput2[18]), .ZN(Red_ToCheckInst_LFInst_52_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_53_LFInst_0_n3), .B(SubCellInput2[22]), .ZN(
        Red_SignaltoCheck[159]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U1 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[21]), .ZN(Red_ToCheckInst_LFInst_53_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_53_LFInst_1_n3), .B(SubCellInput2[23]), .ZN(
        Red_SignaltoCheck[160]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_1_U1 ( .A(SubCellInput2[20]), .B(
        SubCellInput2[21]), .ZN(Red_ToCheckInst_LFInst_53_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_53_LFInst_2_n3), .B(SubCellInput2[23]), .ZN(
        Red_SignaltoCheck[161]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_2_U1 ( .A(SubCellInput2[21]), .B(
        SubCellInput2[22]), .ZN(Red_ToCheckInst_LFInst_53_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_54_LFInst_0_n3), .B(SubCellInput2[26]), .ZN(
        Red_SignaltoCheck[162]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U1 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[25]), .ZN(Red_ToCheckInst_LFInst_54_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_54_LFInst_1_n3), .B(SubCellInput2[27]), .ZN(
        Red_SignaltoCheck[163]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_1_U1 ( .A(SubCellInput2[24]), .B(
        SubCellInput2[25]), .ZN(Red_ToCheckInst_LFInst_54_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_54_LFInst_2_n3), .B(SubCellInput2[27]), .ZN(
        Red_SignaltoCheck[164]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_2_U1 ( .A(SubCellInput2[25]), .B(
        SubCellInput2[26]), .ZN(Red_ToCheckInst_LFInst_54_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_55_LFInst_0_n3), .B(SubCellInput2[30]), .ZN(
        Red_SignaltoCheck[165]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U1 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[29]), .ZN(Red_ToCheckInst_LFInst_55_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_55_LFInst_1_n3), .B(SubCellInput2[31]), .ZN(
        Red_SignaltoCheck[166]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_1_U1 ( .A(SubCellInput2[28]), .B(
        SubCellInput2[29]), .ZN(Red_ToCheckInst_LFInst_55_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_55_LFInst_2_n3), .B(SubCellInput2[31]), .ZN(
        Red_SignaltoCheck[167]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_2_U1 ( .A(SubCellInput2[29]), .B(
        SubCellInput2[30]), .ZN(Red_ToCheckInst_LFInst_55_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_56_LFInst_0_n3), .B(SubCellInput2[34]), .ZN(
        Red_SignaltoCheck[168]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U1 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[33]), .ZN(Red_ToCheckInst_LFInst_56_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_56_LFInst_1_n3), .B(SubCellInput2[35]), .ZN(
        Red_SignaltoCheck[169]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_1_U1 ( .A(SubCellInput2[32]), .B(
        SubCellInput2[33]), .ZN(Red_ToCheckInst_LFInst_56_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_56_LFInst_2_n3), .B(SubCellInput2[35]), .ZN(
        Red_SignaltoCheck[170]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_2_U1 ( .A(SubCellInput2[33]), .B(
        SubCellInput2[34]), .ZN(Red_ToCheckInst_LFInst_56_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_57_LFInst_0_n3), .B(SubCellInput2[38]), .ZN(
        Red_SignaltoCheck[171]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U1 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[37]), .ZN(Red_ToCheckInst_LFInst_57_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_57_LFInst_1_n3), .B(SubCellInput2[39]), .ZN(
        Red_SignaltoCheck[172]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_1_U1 ( .A(SubCellInput2[36]), .B(
        SubCellInput2[37]), .ZN(Red_ToCheckInst_LFInst_57_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_57_LFInst_2_n3), .B(SubCellInput2[39]), .ZN(
        Red_SignaltoCheck[173]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_2_U1 ( .A(SubCellInput2[37]), .B(
        SubCellInput2[38]), .ZN(Red_ToCheckInst_LFInst_57_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_58_LFInst_0_n3), .B(SubCellInput2[42]), .ZN(
        Red_SignaltoCheck[174]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U1 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[41]), .ZN(Red_ToCheckInst_LFInst_58_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_58_LFInst_1_n3), .B(SubCellInput2[43]), .ZN(
        Red_SignaltoCheck[175]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_1_U1 ( .A(SubCellInput2[40]), .B(
        SubCellInput2[41]), .ZN(Red_ToCheckInst_LFInst_58_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_58_LFInst_2_n3), .B(SubCellInput2[43]), .ZN(
        Red_SignaltoCheck[176]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_2_U1 ( .A(SubCellInput2[41]), .B(
        SubCellInput2[42]), .ZN(Red_ToCheckInst_LFInst_58_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_59_LFInst_0_n3), .B(SubCellInput2[46]), .ZN(
        Red_SignaltoCheck[177]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U1 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[45]), .ZN(Red_ToCheckInst_LFInst_59_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_59_LFInst_1_n3), .B(SubCellInput2[47]), .ZN(
        Red_SignaltoCheck[178]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_1_U1 ( .A(SubCellInput2[44]), .B(
        SubCellInput2[45]), .ZN(Red_ToCheckInst_LFInst_59_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_59_LFInst_2_n3), .B(SubCellInput2[47]), .ZN(
        Red_SignaltoCheck[179]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_2_U1 ( .A(SubCellInput2[45]), .B(
        SubCellInput2[46]), .ZN(Red_ToCheckInst_LFInst_59_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_60_LFInst_0_n3), .B(SubCellInput2[50]), .ZN(
        Red_SignaltoCheck[180]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U1 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[49]), .ZN(Red_ToCheckInst_LFInst_60_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_60_LFInst_1_n3), .B(SubCellInput2[51]), .ZN(
        Red_SignaltoCheck[181]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_1_U1 ( .A(SubCellInput2[48]), .B(
        SubCellInput2[49]), .ZN(Red_ToCheckInst_LFInst_60_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_60_LFInst_2_n3), .B(SubCellInput2[51]), .ZN(
        Red_SignaltoCheck[182]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_2_U1 ( .A(SubCellInput2[49]), .B(
        SubCellInput2[50]), .ZN(Red_ToCheckInst_LFInst_60_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_61_LFInst_0_n3), .B(SubCellInput2[54]), .ZN(
        Red_SignaltoCheck[183]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U1 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[53]), .ZN(Red_ToCheckInst_LFInst_61_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_61_LFInst_1_n3), .B(SubCellInput2[55]), .ZN(
        Red_SignaltoCheck[184]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_1_U1 ( .A(SubCellInput2[52]), .B(
        SubCellInput2[53]), .ZN(Red_ToCheckInst_LFInst_61_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_61_LFInst_2_n3), .B(SubCellInput2[55]), .ZN(
        Red_SignaltoCheck[185]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_2_U1 ( .A(SubCellInput2[53]), .B(
        SubCellInput2[54]), .ZN(Red_ToCheckInst_LFInst_61_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_62_LFInst_0_n3), .B(SubCellInput2[58]), .ZN(
        Red_SignaltoCheck[186]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U1 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[57]), .ZN(Red_ToCheckInst_LFInst_62_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_62_LFInst_1_n3), .B(SubCellInput2[59]), .ZN(
        Red_SignaltoCheck[187]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_1_U1 ( .A(SubCellInput2[56]), .B(
        SubCellInput2[57]), .ZN(Red_ToCheckInst_LFInst_62_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_62_LFInst_2_n3), .B(SubCellInput2[59]), .ZN(
        Red_SignaltoCheck[188]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_2_U1 ( .A(SubCellInput2[57]), .B(
        SubCellInput2[58]), .ZN(Red_ToCheckInst_LFInst_62_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_63_LFInst_0_n3), .B(SubCellInput2[62]), .ZN(
        Red_SignaltoCheck[189]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U1 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[61]), .ZN(Red_ToCheckInst_LFInst_63_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_63_LFInst_1_n3), .B(SubCellInput2[63]), .ZN(
        Red_SignaltoCheck[190]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_1_U1 ( .A(SubCellInput2[60]), .B(
        SubCellInput2[61]), .ZN(Red_ToCheckInst_LFInst_63_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_63_LFInst_2_n3), .B(SubCellInput2[63]), .ZN(
        Red_SignaltoCheck[191]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_2_U1 ( .A(SubCellInput2[61]), .B(
        SubCellInput2[62]), .ZN(Red_ToCheckInst_LFInst_63_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_64_LFInst_0_n3), .B(MC_output[2]), .ZN(
        Red_SignaltoCheck[192]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U1 ( .A(MC_output[0]), .B(
        MC_output[1]), .ZN(Red_ToCheckInst_LFInst_64_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_64_LFInst_1_n3), .B(MC_output[3]), .ZN(
        Red_SignaltoCheck[193]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_1_U1 ( .A(MC_output[0]), .B(
        MC_output[1]), .ZN(Red_ToCheckInst_LFInst_64_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_64_LFInst_2_n3), .B(MC_output[3]), .ZN(
        Red_SignaltoCheck[194]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_2_U1 ( .A(MC_output[1]), .B(
        MC_output[2]), .ZN(Red_ToCheckInst_LFInst_64_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_65_LFInst_0_n3), .B(MC_output[6]), .ZN(
        Red_SignaltoCheck[195]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U1 ( .A(MC_output[4]), .B(
        MC_output[5]), .ZN(Red_ToCheckInst_LFInst_65_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_65_LFInst_1_n3), .B(MC_output[7]), .ZN(
        Red_SignaltoCheck[196]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_1_U1 ( .A(MC_output[4]), .B(
        MC_output[5]), .ZN(Red_ToCheckInst_LFInst_65_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_65_LFInst_2_n3), .B(MC_output[7]), .ZN(
        Red_SignaltoCheck[197]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_2_U1 ( .A(MC_output[5]), .B(
        MC_output[6]), .ZN(Red_ToCheckInst_LFInst_65_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_66_LFInst_0_n3), .B(MC_output[10]), .ZN(
        Red_SignaltoCheck[198]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U1 ( .A(MC_output[8]), .B(
        MC_output[9]), .ZN(Red_ToCheckInst_LFInst_66_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_66_LFInst_1_n3), .B(MC_output[11]), .ZN(
        Red_SignaltoCheck[199]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_1_U1 ( .A(MC_output[8]), .B(
        MC_output[9]), .ZN(Red_ToCheckInst_LFInst_66_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_66_LFInst_2_n3), .B(MC_output[11]), .ZN(
        Red_SignaltoCheck[200]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_2_U1 ( .A(MC_output[9]), .B(
        MC_output[10]), .ZN(Red_ToCheckInst_LFInst_66_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_67_LFInst_0_n3), .B(MC_output[14]), .ZN(
        Red_SignaltoCheck[201]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U1 ( .A(MC_output[12]), .B(
        MC_output[13]), .ZN(Red_ToCheckInst_LFInst_67_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_67_LFInst_1_n3), .B(MC_output[15]), .ZN(
        Red_SignaltoCheck[202]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_1_U1 ( .A(MC_output[12]), .B(
        MC_output[13]), .ZN(Red_ToCheckInst_LFInst_67_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_67_LFInst_2_n3), .B(MC_output[15]), .ZN(
        Red_SignaltoCheck[203]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_2_U1 ( .A(MC_output[13]), .B(
        MC_output[14]), .ZN(Red_ToCheckInst_LFInst_67_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_68_LFInst_0_n3), .B(MC_output[18]), .ZN(
        Red_SignaltoCheck[204]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U1 ( .A(MC_output[16]), .B(
        MC_output[17]), .ZN(Red_ToCheckInst_LFInst_68_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_68_LFInst_1_n3), .B(MC_output[19]), .ZN(
        Red_SignaltoCheck[205]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_1_U1 ( .A(MC_output[16]), .B(
        MC_output[17]), .ZN(Red_ToCheckInst_LFInst_68_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_68_LFInst_2_n3), .B(MC_output[19]), .ZN(
        Red_SignaltoCheck[206]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_2_U1 ( .A(MC_output[17]), .B(
        MC_output[18]), .ZN(Red_ToCheckInst_LFInst_68_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_69_LFInst_0_n3), .B(MC_output[22]), .ZN(
        Red_SignaltoCheck[207]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U1 ( .A(MC_output[20]), .B(
        MC_output[21]), .ZN(Red_ToCheckInst_LFInst_69_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_69_LFInst_1_n3), .B(MC_output[23]), .ZN(
        Red_SignaltoCheck[208]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_1_U1 ( .A(MC_output[20]), .B(
        MC_output[21]), .ZN(Red_ToCheckInst_LFInst_69_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_69_LFInst_2_n3), .B(MC_output[23]), .ZN(
        Red_SignaltoCheck[209]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_2_U1 ( .A(MC_output[21]), .B(
        MC_output[22]), .ZN(Red_ToCheckInst_LFInst_69_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_70_LFInst_0_n3), .B(MC_output[26]), .ZN(
        Red_SignaltoCheck[210]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U1 ( .A(MC_output[24]), .B(
        MC_output[25]), .ZN(Red_ToCheckInst_LFInst_70_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_70_LFInst_1_n3), .B(MC_output[27]), .ZN(
        Red_SignaltoCheck[211]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_1_U1 ( .A(MC_output[24]), .B(
        MC_output[25]), .ZN(Red_ToCheckInst_LFInst_70_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_70_LFInst_2_n3), .B(MC_output[27]), .ZN(
        Red_SignaltoCheck[212]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_2_U1 ( .A(MC_output[25]), .B(
        MC_output[26]), .ZN(Red_ToCheckInst_LFInst_70_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_71_LFInst_0_n3), .B(MC_output[30]), .ZN(
        Red_SignaltoCheck[213]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U1 ( .A(MC_output[28]), .B(
        MC_output[29]), .ZN(Red_ToCheckInst_LFInst_71_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_71_LFInst_1_n3), .B(MC_output[31]), .ZN(
        Red_SignaltoCheck[214]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_1_U1 ( .A(MC_output[28]), .B(
        MC_output[29]), .ZN(Red_ToCheckInst_LFInst_71_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_71_LFInst_2_n3), .B(MC_output[31]), .ZN(
        Red_SignaltoCheck[215]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_2_U1 ( .A(MC_output[29]), .B(
        MC_output[30]), .ZN(Red_ToCheckInst_LFInst_71_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_72_LFInst_0_n3), .B(MC_output[34]), .ZN(
        Red_SignaltoCheck[216]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U1 ( .A(MC_output[32]), .B(
        MC_output[33]), .ZN(Red_ToCheckInst_LFInst_72_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_72_LFInst_1_n3), .B(MC_output[35]), .ZN(
        Red_SignaltoCheck[217]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_1_U1 ( .A(MC_output[32]), .B(
        MC_output[33]), .ZN(Red_ToCheckInst_LFInst_72_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_72_LFInst_2_n3), .B(MC_output[35]), .ZN(
        Red_SignaltoCheck[218]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_2_U1 ( .A(MC_output[33]), .B(
        MC_output[34]), .ZN(Red_ToCheckInst_LFInst_72_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_73_LFInst_0_n3), .B(MC_output[38]), .ZN(
        Red_SignaltoCheck[219]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U1 ( .A(MC_output[36]), .B(
        MC_output[37]), .ZN(Red_ToCheckInst_LFInst_73_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_73_LFInst_1_n3), .B(MC_output[39]), .ZN(
        Red_SignaltoCheck[220]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_1_U1 ( .A(MC_output[36]), .B(
        MC_output[37]), .ZN(Red_ToCheckInst_LFInst_73_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_73_LFInst_2_n3), .B(MC_output[39]), .ZN(
        Red_SignaltoCheck[221]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_2_U1 ( .A(MC_output[37]), .B(
        MC_output[38]), .ZN(Red_ToCheckInst_LFInst_73_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_74_LFInst_0_n3), .B(MC_output[42]), .ZN(
        Red_SignaltoCheck[222]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U1 ( .A(MC_output[40]), .B(
        MC_output[41]), .ZN(Red_ToCheckInst_LFInst_74_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_74_LFInst_1_n3), .B(MC_output[43]), .ZN(
        Red_SignaltoCheck[223]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_1_U1 ( .A(MC_output[40]), .B(
        MC_output[41]), .ZN(Red_ToCheckInst_LFInst_74_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_74_LFInst_2_n3), .B(MC_output[43]), .ZN(
        Red_SignaltoCheck[224]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_2_U1 ( .A(MC_output[41]), .B(
        MC_output[42]), .ZN(Red_ToCheckInst_LFInst_74_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_75_LFInst_0_n3), .B(MC_output[46]), .ZN(
        Red_SignaltoCheck[225]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U1 ( .A(MC_output[44]), .B(
        MC_output[45]), .ZN(Red_ToCheckInst_LFInst_75_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_75_LFInst_1_n3), .B(MC_output[47]), .ZN(
        Red_SignaltoCheck[226]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_1_U1 ( .A(MC_output[44]), .B(
        MC_output[45]), .ZN(Red_ToCheckInst_LFInst_75_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_75_LFInst_2_n3), .B(MC_output[47]), .ZN(
        Red_SignaltoCheck[227]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_2_U1 ( .A(MC_output[45]), .B(
        MC_output[46]), .ZN(Red_ToCheckInst_LFInst_75_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_76_LFInst_0_n3), .B(MC_output[50]), .ZN(
        Red_SignaltoCheck[228]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U1 ( .A(MC_output[48]), .B(
        MC_output[49]), .ZN(Red_ToCheckInst_LFInst_76_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_76_LFInst_1_n3), .B(MC_output[51]), .ZN(
        Red_SignaltoCheck[229]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_1_U1 ( .A(MC_output[48]), .B(
        MC_output[49]), .ZN(Red_ToCheckInst_LFInst_76_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_76_LFInst_2_n3), .B(MC_output[51]), .ZN(
        Red_SignaltoCheck[230]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_2_U1 ( .A(MC_output[49]), .B(
        MC_output[50]), .ZN(Red_ToCheckInst_LFInst_76_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_77_LFInst_0_n3), .B(MC_output[54]), .ZN(
        Red_SignaltoCheck[231]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U1 ( .A(MC_output[52]), .B(
        MC_output[53]), .ZN(Red_ToCheckInst_LFInst_77_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_77_LFInst_1_n3), .B(MC_output[55]), .ZN(
        Red_SignaltoCheck[232]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_1_U1 ( .A(MC_output[52]), .B(
        MC_output[53]), .ZN(Red_ToCheckInst_LFInst_77_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_77_LFInst_2_n3), .B(MC_output[55]), .ZN(
        Red_SignaltoCheck[233]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_2_U1 ( .A(MC_output[53]), .B(
        MC_output[54]), .ZN(Red_ToCheckInst_LFInst_77_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_78_LFInst_0_n3), .B(MC_output[58]), .ZN(
        Red_SignaltoCheck[234]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U1 ( .A(MC_output[56]), .B(
        MC_output[57]), .ZN(Red_ToCheckInst_LFInst_78_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_78_LFInst_1_n3), .B(MC_output[59]), .ZN(
        Red_SignaltoCheck[235]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_1_U1 ( .A(MC_output[56]), .B(
        MC_output[57]), .ZN(Red_ToCheckInst_LFInst_78_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_78_LFInst_2_n3), .B(MC_output[59]), .ZN(
        Red_SignaltoCheck[236]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_2_U1 ( .A(MC_output[57]), .B(
        MC_output[58]), .ZN(Red_ToCheckInst_LFInst_78_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_79_LFInst_0_n3), .B(MC_output[62]), .ZN(
        Red_SignaltoCheck[237]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U1 ( .A(MC_output[60]), .B(
        MC_output[61]), .ZN(Red_ToCheckInst_LFInst_79_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_79_LFInst_1_n3), .B(MC_output[63]), .ZN(
        Red_SignaltoCheck[238]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_1_U1 ( .A(MC_output[60]), .B(
        MC_output[61]), .ZN(Red_ToCheckInst_LFInst_79_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_79_LFInst_2_n3), .B(MC_output[63]), .ZN(
        Red_SignaltoCheck[239]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_2_U1 ( .A(MC_output[61]), .B(
        MC_output[62]), .ZN(Red_ToCheckInst_LFInst_79_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_80_LFInst_0_n3), .B(MCInst_MC3_v3_0[3]), .ZN(
        Red_SignaltoCheck[240]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_80_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_80_LFInst_1_n3), .B(Red_MCInst_MC3_v3_1[2]), 
        .ZN(Red_SignaltoCheck[241]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_1_U1 ( .A(MCInst_MC3_v3_2[3]), .B(
        Red_MCInst_MC3_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_80_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_80_LFInst_2_n3), .B(Red_MCInst_MC3_v3_1[2]), 
        .ZN(Red_SignaltoCheck[242]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_2_U1 ( .A(Red_MCInst_MC3_v3_3[2]), 
        .B(MCInst_MC3_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_80_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_81_LFInst_0_n3), .B(MCInst_MC2_v3_0[3]), .ZN(
        Red_SignaltoCheck[243]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_81_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_81_LFInst_1_n3), .B(Red_MCInst_MC2_v3_1[2]), 
        .ZN(Red_SignaltoCheck[244]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_1_U1 ( .A(MCInst_MC2_v3_2[3]), .B(
        Red_MCInst_MC2_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_81_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_81_LFInst_2_n3), .B(Red_MCInst_MC2_v3_1[2]), 
        .ZN(Red_SignaltoCheck[245]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_2_U1 ( .A(Red_MCInst_MC2_v3_3[2]), 
        .B(MCInst_MC2_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_81_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_82_LFInst_0_n3), .B(MCInst_MC1_v3_0[3]), .ZN(
        Red_SignaltoCheck[246]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_82_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_82_LFInst_1_n3), .B(Red_MCInst_MC1_v3_1[2]), 
        .ZN(Red_SignaltoCheck[247]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_1_U1 ( .A(MCInst_MC1_v3_2[3]), .B(
        Red_MCInst_MC1_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_82_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_82_LFInst_2_n3), .B(Red_MCInst_MC1_v3_1[2]), 
        .ZN(Red_SignaltoCheck[248]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_2_U1 ( .A(Red_MCInst_MC1_v3_3[2]), 
        .B(MCInst_MC1_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_82_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_83_LFInst_0_n3), .B(MCInst_MC0_v3_0[3]), .ZN(
        Red_SignaltoCheck[249]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_83_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_83_LFInst_1_n3), .B(Red_MCInst_MC0_v3_1[2]), 
        .ZN(Red_SignaltoCheck[250]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_1_U1 ( .A(MCInst_MC0_v3_2[3]), .B(
        Red_MCInst_MC0_v3_3[2]), .ZN(Red_ToCheckInst_LFInst_83_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_83_LFInst_2_n3), .B(Red_MCInst_MC0_v3_1[2]), 
        .ZN(Red_SignaltoCheck[251]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_2_U1 ( .A(Red_MCInst_MC0_v3_3[2]), 
        .B(MCInst_MC0_v3_0[3]), .ZN(Red_ToCheckInst_LFInst_83_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_84_LFInst_0_n3), .B(MCInst_MC3_v2_0[3]), .ZN(
        Red_SignaltoCheck[252]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U1 ( .A(ShiftRowsOutput[16]), 
        .B(MCInst_MC3_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_84_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_84_LFInst_1_n3), .B(Red_MCInst_MC3_v2_2[1]), 
        .ZN(Red_SignaltoCheck[253]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_1_U1 ( .A(ShiftRowsOutput[16]), 
        .B(MCInst_MC3_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_84_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_84_LFInst_2_n3), .B(Red_MCInst_MC3_v2_2[1]), 
        .ZN(Red_SignaltoCheck[254]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_2_U1 ( .A(MCInst_MC3_v2_0[2]), .B(
        MCInst_MC3_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_84_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_85_LFInst_0_n3), .B(MCInst_MC2_v2_0[3]), .ZN(
        Red_SignaltoCheck[255]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U1 ( .A(ShiftRowsOutput[20]), 
        .B(MCInst_MC2_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_85_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_85_LFInst_1_n3), .B(Red_MCInst_MC2_v2_2[1]), 
        .ZN(Red_SignaltoCheck[256]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_1_U1 ( .A(ShiftRowsOutput[20]), 
        .B(MCInst_MC2_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_85_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_85_LFInst_2_n3), .B(Red_MCInst_MC2_v2_2[1]), 
        .ZN(Red_SignaltoCheck[257]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_2_U1 ( .A(MCInst_MC2_v2_0[2]), .B(
        MCInst_MC2_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_85_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_86_LFInst_0_n3), .B(MCInst_MC1_v2_0[3]), .ZN(
        Red_SignaltoCheck[258]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U1 ( .A(ShiftRowsOutput[24]), 
        .B(MCInst_MC1_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_86_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_86_LFInst_1_n3), .B(Red_MCInst_MC1_v2_2[1]), 
        .ZN(Red_SignaltoCheck[259]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_1_U1 ( .A(ShiftRowsOutput[24]), 
        .B(MCInst_MC1_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_86_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_86_LFInst_2_n3), .B(Red_MCInst_MC1_v2_2[1]), 
        .ZN(Red_SignaltoCheck[260]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_2_U1 ( .A(MCInst_MC1_v2_0[2]), .B(
        MCInst_MC1_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_86_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_87_LFInst_0_n3), .B(MCInst_MC0_v2_0[3]), .ZN(
        Red_SignaltoCheck[261]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U1 ( .A(ShiftRowsOutput[28]), 
        .B(MCInst_MC0_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_87_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_87_LFInst_1_n3), .B(Red_MCInst_MC0_v2_2[1]), 
        .ZN(Red_SignaltoCheck[262]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_1_U1 ( .A(ShiftRowsOutput[28]), 
        .B(MCInst_MC0_v2_0[2]), .ZN(Red_ToCheckInst_LFInst_87_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_87_LFInst_2_n3), .B(Red_MCInst_MC0_v2_2[1]), 
        .ZN(Red_SignaltoCheck[263]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_2_U1 ( .A(MCInst_MC0_v2_0[2]), .B(
        MCInst_MC0_v2_0[3]), .ZN(Red_ToCheckInst_LFInst_87_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_88_LFInst_0_n3), .B(MCInst_MC3_v1_3[3]), .ZN(
        Red_SignaltoCheck[264]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_88_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_88_LFInst_1_n3), .B(Red_MCInst_MC3_v1_1[2]), 
        .ZN(Red_SignaltoCheck[265]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_1_U1 ( .A(MCInst_MC3_v1_0_0_), .B(
        MCInst_MC3_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_88_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_88_LFInst_2_n3), .B(Red_MCInst_MC3_v1_1[2]), 
        .ZN(Red_SignaltoCheck[266]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_2_U1 ( .A(MCInst_MC3_v1_3[2]), .B(
        MCInst_MC3_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_88_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_89_LFInst_0_n3), .B(MCInst_MC2_v1_3[3]), .ZN(
        Red_SignaltoCheck[267]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_89_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_89_LFInst_1_n3), .B(Red_MCInst_MC2_v1_1[2]), 
        .ZN(Red_SignaltoCheck[268]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_1_U1 ( .A(MCInst_MC2_v1_0_0_), .B(
        MCInst_MC2_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_89_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_89_LFInst_2_n3), .B(Red_MCInst_MC2_v1_1[2]), 
        .ZN(Red_SignaltoCheck[269]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_2_U1 ( .A(MCInst_MC2_v1_3[2]), .B(
        MCInst_MC2_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_89_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_90_LFInst_0_n3), .B(MCInst_MC1_v1_3[3]), .ZN(
        Red_SignaltoCheck[270]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_90_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_90_LFInst_1_n3), .B(Red_MCInst_MC1_v1_1[2]), 
        .ZN(Red_SignaltoCheck[271]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_1_U1 ( .A(MCInst_MC1_v1_0_0_), .B(
        MCInst_MC1_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_90_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_90_LFInst_2_n3), .B(Red_MCInst_MC1_v1_1[2]), 
        .ZN(Red_SignaltoCheck[272]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_2_U1 ( .A(MCInst_MC1_v1_3[2]), .B(
        MCInst_MC1_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_90_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_91_LFInst_0_n3), .B(MCInst_MC0_v1_3[3]), .ZN(
        Red_SignaltoCheck[273]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_91_LFInst_0_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_91_LFInst_1_n3), .B(Red_MCInst_MC0_v1_1[2]), 
        .ZN(Red_SignaltoCheck[274]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_1_U1 ( .A(MCInst_MC0_v1_0_0_), .B(
        MCInst_MC0_v1_3[2]), .ZN(Red_ToCheckInst_LFInst_91_LFInst_1_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_91_LFInst_2_n3), .B(Red_MCInst_MC0_v1_1[2]), 
        .ZN(Red_SignaltoCheck[275]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_2_U1 ( .A(MCInst_MC0_v1_3[2]), .B(
        MCInst_MC0_v1_3[3]), .ZN(Red_ToCheckInst_LFInst_91_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_92_LFInst_0_n3), .B(MCInst_MC3_v0_3[3]), .ZN(
        Red_SignaltoCheck[276]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U1 ( .A(Red_MCInst_MC3_v0_0[0]), 
        .B(Red_MCInst_MC3_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_92_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_92_LFInst_1_n3), .B(Red_MCInst_MC3_v0_1[0]), 
        .ZN(Red_SignaltoCheck[277]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_1_U1 ( .A(Red_MCInst_MC3_v0_0[0]), 
        .B(Red_MCInst_MC3_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_92_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_92_LFInst_2_n3), .B(Red_MCInst_MC3_v0_1[0]), 
        .ZN(Red_SignaltoCheck[278]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_2_U1 ( .A(Red_MCInst_MC3_v0_2[2]), 
        .B(MCInst_MC3_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_92_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_93_LFInst_0_n3), .B(MCInst_MC2_v0_3[3]), .ZN(
        Red_SignaltoCheck[279]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U1 ( .A(Red_MCInst_MC2_v0_0[0]), 
        .B(Red_MCInst_MC2_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_93_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_93_LFInst_1_n3), .B(Red_MCInst_MC2_v0_1[0]), 
        .ZN(Red_SignaltoCheck[280]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_1_U1 ( .A(Red_MCInst_MC2_v0_0[0]), 
        .B(Red_MCInst_MC2_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_93_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_93_LFInst_2_n3), .B(Red_MCInst_MC2_v0_1[0]), 
        .ZN(Red_SignaltoCheck[281]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_2_U1 ( .A(Red_MCInst_MC2_v0_2[2]), 
        .B(MCInst_MC2_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_93_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_94_LFInst_0_n3), .B(MCInst_MC1_v0_3[3]), .ZN(
        Red_SignaltoCheck[282]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U1 ( .A(Red_MCInst_MC1_v0_0[0]), 
        .B(Red_MCInst_MC1_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_94_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_94_LFInst_1_n3), .B(Red_MCInst_MC1_v0_1[0]), 
        .ZN(Red_SignaltoCheck[283]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_1_U1 ( .A(Red_MCInst_MC1_v0_0[0]), 
        .B(Red_MCInst_MC1_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_94_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_94_LFInst_2_n3), .B(Red_MCInst_MC1_v0_1[0]), 
        .ZN(Red_SignaltoCheck[284]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_2_U1 ( .A(Red_MCInst_MC1_v0_2[2]), 
        .B(MCInst_MC1_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_94_LFInst_2_n3) );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_95_LFInst_0_n3), .B(MCInst_MC0_v0_3[3]), .ZN(
        Red_SignaltoCheck[285]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U1 ( .A(Red_MCInst_MC0_v0_0[0]), 
        .B(Red_MCInst_MC0_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_95_LFInst_0_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_95_LFInst_1_n3), .B(Red_MCInst_MC0_v0_1[0]), 
        .ZN(Red_SignaltoCheck[286]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_1_U1 ( .A(Red_MCInst_MC0_v0_0[0]), 
        .B(Red_MCInst_MC0_v0_2[2]), .ZN(Red_ToCheckInst_LFInst_95_LFInst_1_n3)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_95_LFInst_2_n3), .B(Red_MCInst_MC0_v0_1[0]), 
        .ZN(Red_SignaltoCheck[287]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_2_U1 ( .A(Red_MCInst_MC0_v0_2[2]), 
        .B(MCInst_MC0_v0_3[3]), .ZN(Red_ToCheckInst_LFInst_95_LFInst_2_n3) );
  NOR2_X1 Check1_CheckInst_0_U191 ( .A1(Check1_CheckInst_0_n190), .A2(
        Check1_CheckInst_0_n189), .ZN(Error[0]) );
  NAND2_X1 Check1_CheckInst_0_U190 ( .A1(Check1_CheckInst_0_n188), .A2(
        Check1_CheckInst_0_n187), .ZN(Check1_CheckInst_0_n189) );
  NOR2_X1 Check1_CheckInst_0_U189 ( .A1(Check1_CheckInst_0_n186), .A2(
        Check1_CheckInst_0_n185), .ZN(Check1_CheckInst_0_n187) );
  NAND2_X1 Check1_CheckInst_0_U188 ( .A1(Check1_CheckInst_0_n184), .A2(
        Check1_CheckInst_0_n183), .ZN(Check1_CheckInst_0_n185) );
  NOR2_X1 Check1_CheckInst_0_U187 ( .A1(Check1_CheckInst_0_n182), .A2(
        Check1_CheckInst_0_n181), .ZN(Check1_CheckInst_0_n183) );
  NAND2_X1 Check1_CheckInst_0_U186 ( .A1(Check1_CheckInst_0_n180), .A2(
        Check1_CheckInst_0_n179), .ZN(Check1_CheckInst_0_n181) );
  NOR2_X1 Check1_CheckInst_0_U185 ( .A1(Check1_CheckInst_0_n178), .A2(
        Check1_CheckInst_0_n177), .ZN(Check1_CheckInst_0_n179) );
  NAND2_X1 Check1_CheckInst_0_U184 ( .A1(Check1_CheckInst_0_n176), .A2(
        Check1_CheckInst_0_n175), .ZN(Check1_CheckInst_0_n177) );
  NOR2_X1 Check1_CheckInst_0_U183 ( .A1(Check1_CheckInst_0_n174), .A2(
        Check1_CheckInst_0_n173), .ZN(Check1_CheckInst_0_n175) );
  NAND2_X1 Check1_CheckInst_0_U182 ( .A1(Check1_CheckInst_0_n172), .A2(
        Check1_CheckInst_0_n171), .ZN(Check1_CheckInst_0_n173) );
  XNOR2_X1 Check1_CheckInst_0_U181 ( .A(Red_ShiftRowsOutput[30]), .B(
        Red_SignaltoCheck[270]), .ZN(Check1_CheckInst_0_n171) );
  XNOR2_X1 Check1_CheckInst_0_U180 ( .A(Red_ShiftRowsOutput[36]), .B(
        Red_SignaltoCheck[276]), .ZN(Check1_CheckInst_0_n172) );
  NAND2_X1 Check1_CheckInst_0_U179 ( .A1(Check1_CheckInst_0_n170), .A2(
        Check1_CheckInst_0_n169), .ZN(Check1_CheckInst_0_n174) );
  XNOR2_X1 Check1_CheckInst_0_U178 ( .A(Red_ShiftRowsOutput[27]), .B(
        Red_SignaltoCheck[267]), .ZN(Check1_CheckInst_0_n169) );
  XNOR2_X1 Check1_CheckInst_0_U177 ( .A(Red_ShiftRowsOutput[33]), .B(
        Red_SignaltoCheck[273]), .ZN(Check1_CheckInst_0_n170) );
  NOR2_X1 Check1_CheckInst_0_U176 ( .A1(Check1_CheckInst_0_n168), .A2(
        Check1_CheckInst_0_n167), .ZN(Check1_CheckInst_0_n176) );
  XOR2_X1 Check1_CheckInst_0_U175 ( .A(Red_MC_output[36]), .B(
        Red_SignaltoCheck[228]), .Z(Check1_CheckInst_0_n167) );
  XOR2_X1 Check1_CheckInst_0_U174 ( .A(Red_MC_output[33]), .B(
        Red_SignaltoCheck[225]), .Z(Check1_CheckInst_0_n168) );
  NAND2_X1 Check1_CheckInst_0_U173 ( .A1(Check1_CheckInst_0_n166), .A2(
        Check1_CheckInst_0_n165), .ZN(Check1_CheckInst_0_n178) );
  XNOR2_X1 Check1_CheckInst_0_U172 ( .A(Red_MC_output[24]), .B(
        Red_SignaltoCheck[216]), .ZN(Check1_CheckInst_0_n165) );
  XNOR2_X1 Check1_CheckInst_0_U171 ( .A(Red_MC_output[30]), .B(
        Red_SignaltoCheck[222]), .ZN(Check1_CheckInst_0_n166) );
  NOR2_X1 Check1_CheckInst_0_U170 ( .A1(Check1_CheckInst_0_n164), .A2(
        Check1_CheckInst_0_n163), .ZN(Check1_CheckInst_0_n180) );
  NAND2_X1 Check1_CheckInst_0_U169 ( .A1(Check1_CheckInst_0_n162), .A2(
        Check1_CheckInst_0_n161), .ZN(Check1_CheckInst_0_n163) );
  NOR2_X1 Check1_CheckInst_0_U168 ( .A1(Check1_CheckInst_0_n160), .A2(
        Check1_CheckInst_0_n159), .ZN(Check1_CheckInst_0_n161) );
  NAND2_X1 Check1_CheckInst_0_U167 ( .A1(Check1_CheckInst_0_n158), .A2(
        Check1_CheckInst_0_n157), .ZN(Check1_CheckInst_0_n159) );
  XNOR2_X1 Check1_CheckInst_0_U166 ( .A(Red_MC_output[21]), .B(
        Red_SignaltoCheck[213]), .ZN(Check1_CheckInst_0_n157) );
  XNOR2_X1 Check1_CheckInst_0_U165 ( .A(Red_MC_output[27]), .B(
        Red_SignaltoCheck[219]), .ZN(Check1_CheckInst_0_n158) );
  NAND2_X1 Check1_CheckInst_0_U164 ( .A1(Check1_CheckInst_0_n156), .A2(
        Check1_CheckInst_0_n155), .ZN(Check1_CheckInst_0_n160) );
  XNOR2_X1 Check1_CheckInst_0_U163 ( .A(Red_ShiftRowsOutput[6]), .B(
        Red_SignaltoCheck[246]), .ZN(Check1_CheckInst_0_n155) );
  XNOR2_X1 Check1_CheckInst_0_U162 ( .A(Red_ShiftRowsOutput[3]), .B(
        Red_SignaltoCheck[243]), .ZN(Check1_CheckInst_0_n156) );
  NOR2_X1 Check1_CheckInst_0_U161 ( .A1(Check1_CheckInst_0_n154), .A2(
        Check1_CheckInst_0_n153), .ZN(Check1_CheckInst_0_n162) );
  XOR2_X1 Check1_CheckInst_0_U160 ( .A(Red_MC_output[42]), .B(
        Red_SignaltoCheck[234]), .Z(Check1_CheckInst_0_n153) );
  XOR2_X1 Check1_CheckInst_0_U159 ( .A(Red_ShiftRowsOutput[0]), .B(
        Red_SignaltoCheck[240]), .Z(Check1_CheckInst_0_n154) );
  NAND2_X1 Check1_CheckInst_0_U158 ( .A1(Check1_CheckInst_0_n152), .A2(
        Check1_CheckInst_0_n151), .ZN(Check1_CheckInst_0_n164) );
  XNOR2_X1 Check1_CheckInst_0_U157 ( .A(Red_MC_output[39]), .B(
        Red_SignaltoCheck[231]), .ZN(Check1_CheckInst_0_n151) );
  XNOR2_X1 Check1_CheckInst_0_U156 ( .A(Red_MC_output[45]), .B(
        Red_SignaltoCheck[237]), .ZN(Check1_CheckInst_0_n152) );
  NAND2_X1 Check1_CheckInst_0_U155 ( .A1(Check1_CheckInst_0_n150), .A2(
        Check1_CheckInst_0_n149), .ZN(Check1_CheckInst_0_n182) );
  NOR2_X1 Check1_CheckInst_0_U154 ( .A1(Check1_CheckInst_0_n148), .A2(
        Check1_CheckInst_0_n147), .ZN(Check1_CheckInst_0_n149) );
  NAND2_X1 Check1_CheckInst_0_U153 ( .A1(Check1_CheckInst_0_n146), .A2(
        Check1_CheckInst_0_n145), .ZN(Check1_CheckInst_0_n147) );
  NOR2_X1 Check1_CheckInst_0_U152 ( .A1(Check1_CheckInst_0_n144), .A2(
        Check1_CheckInst_0_n143), .ZN(Check1_CheckInst_0_n145) );
  XOR2_X1 Check1_CheckInst_0_U151 ( .A(Red_MC_output2[45]), .B(
        Red_SignaltoCheck[93]), .Z(Check1_CheckInst_0_n143) );
  XOR2_X1 Check1_CheckInst_0_U150 ( .A(Red_MC_output2[42]), .B(
        Red_SignaltoCheck[90]), .Z(Check1_CheckInst_0_n144) );
  NOR2_X1 Check1_CheckInst_0_U149 ( .A1(Check1_CheckInst_0_n142), .A2(
        Check1_CheckInst_0_n141), .ZN(Check1_CheckInst_0_n146) );
  XOR2_X1 Check1_CheckInst_0_U148 ( .A(Red_ShiftRowsOutput2[3]), .B(
        Red_SignaltoCheck[99]), .Z(Check1_CheckInst_0_n141) );
  XOR2_X1 Check1_CheckInst_0_U147 ( .A(Red_MC_output2[39]), .B(
        Red_SignaltoCheck[87]), .Z(Check1_CheckInst_0_n142) );
  NAND2_X1 Check1_CheckInst_0_U146 ( .A1(Check1_CheckInst_0_n140), .A2(
        Check1_CheckInst_0_n139), .ZN(Check1_CheckInst_0_n148) );
  XNOR2_X1 Check1_CheckInst_0_U145 ( .A(Red_ShiftRowsOutput2[0]), .B(
        Red_SignaltoCheck[96]), .ZN(Check1_CheckInst_0_n139) );
  XNOR2_X1 Check1_CheckInst_0_U144 ( .A(Red_ShiftRowsOutput2[6]), .B(
        Red_SignaltoCheck[102]), .ZN(Check1_CheckInst_0_n140) );
  NOR2_X1 Check1_CheckInst_0_U143 ( .A1(Check1_CheckInst_0_n138), .A2(
        Check1_CheckInst_0_n137), .ZN(Check1_CheckInst_0_n150) );
  XOR2_X1 Check1_CheckInst_0_U142 ( .A(Red_MC_output2[27]), .B(
        Red_SignaltoCheck[75]), .Z(Check1_CheckInst_0_n137) );
  XOR2_X1 Check1_CheckInst_0_U141 ( .A(Red_MC_output2[24]), .B(
        Red_SignaltoCheck[72]), .Z(Check1_CheckInst_0_n138) );
  NOR2_X1 Check1_CheckInst_0_U140 ( .A1(Check1_CheckInst_0_n136), .A2(
        Check1_CheckInst_0_n135), .ZN(Check1_CheckInst_0_n184) );
  NAND2_X1 Check1_CheckInst_0_U139 ( .A1(Check1_CheckInst_0_n134), .A2(
        Check1_CheckInst_0_n133), .ZN(Check1_CheckInst_0_n135) );
  NOR2_X1 Check1_CheckInst_0_U138 ( .A1(Check1_CheckInst_0_n132), .A2(
        Check1_CheckInst_0_n131), .ZN(Check1_CheckInst_0_n133) );
  NAND2_X1 Check1_CheckInst_0_U137 ( .A1(Check1_CheckInst_0_n130), .A2(
        Check1_CheckInst_0_n129), .ZN(Check1_CheckInst_0_n131) );
  XNOR2_X1 Check1_CheckInst_0_U136 ( .A(Red_MC_output2[33]), .B(
        Red_SignaltoCheck[81]), .ZN(Check1_CheckInst_0_n129) );
  XNOR2_X1 Check1_CheckInst_0_U135 ( .A(Red_MC_output2[21]), .B(
        Red_SignaltoCheck[69]), .ZN(Check1_CheckInst_0_n130) );
  NAND2_X1 Check1_CheckInst_0_U134 ( .A1(Check1_CheckInst_0_n128), .A2(
        Check1_CheckInst_0_n127), .ZN(Check1_CheckInst_0_n132) );
  XNOR2_X1 Check1_CheckInst_0_U133 ( .A(Red_MC_output2[30]), .B(
        Red_SignaltoCheck[78]), .ZN(Check1_CheckInst_0_n127) );
  XNOR2_X1 Check1_CheckInst_0_U132 ( .A(Red_MC_output2[36]), .B(
        Red_SignaltoCheck[84]), .ZN(Check1_CheckInst_0_n128) );
  NOR2_X1 Check1_CheckInst_0_U131 ( .A1(Check1_CheckInst_0_n126), .A2(
        Check1_CheckInst_0_n125), .ZN(Check1_CheckInst_0_n134) );
  XOR2_X1 Check1_CheckInst_0_U130 ( .A(Red_ShiftRowsOutput2[33]), .B(
        Red_SignaltoCheck[129]), .Z(Check1_CheckInst_0_n125) );
  XOR2_X1 Check1_CheckInst_0_U129 ( .A(Red_ShiftRowsOutput2[30]), .B(
        Red_SignaltoCheck[126]), .Z(Check1_CheckInst_0_n126) );
  NAND2_X1 Check1_CheckInst_0_U128 ( .A1(Check1_CheckInst_0_n124), .A2(
        Check1_CheckInst_0_n123), .ZN(Check1_CheckInst_0_n136) );
  XNOR2_X1 Check1_CheckInst_0_U127 ( .A(Red_ShiftRowsOutput2[39]), .B(
        Red_SignaltoCheck[135]), .ZN(Check1_CheckInst_0_n123) );
  XNOR2_X1 Check1_CheckInst_0_U126 ( .A(Red_ShiftRowsOutput2[27]), .B(
        Red_SignaltoCheck[123]), .ZN(Check1_CheckInst_0_n124) );
  NAND2_X1 Check1_CheckInst_0_U125 ( .A1(Check1_CheckInst_0_n122), .A2(
        Check1_CheckInst_0_n121), .ZN(Check1_CheckInst_0_n186) );
  NOR2_X1 Check1_CheckInst_0_U124 ( .A1(Check1_CheckInst_0_n120), .A2(
        Check1_CheckInst_0_n119), .ZN(Check1_CheckInst_0_n121) );
  NAND2_X1 Check1_CheckInst_0_U123 ( .A1(Check1_CheckInst_0_n118), .A2(
        Check1_CheckInst_0_n117), .ZN(Check1_CheckInst_0_n119) );
  NOR2_X1 Check1_CheckInst_0_U122 ( .A1(Check1_CheckInst_0_n116), .A2(
        Check1_CheckInst_0_n115), .ZN(Check1_CheckInst_0_n117) );
  XOR2_X1 Check1_CheckInst_0_U121 ( .A(Red_SubCellInput2[12]), .B(
        Red_SignaltoCheck[156]), .Z(Check1_CheckInst_0_n115) );
  XOR2_X1 Check1_CheckInst_0_U120 ( .A(Red_SubCellInput2[9]), .B(
        Red_SignaltoCheck[153]), .Z(Check1_CheckInst_0_n116) );
  XNOR2_X1 Check1_CheckInst_0_U119 ( .A(Red_SubCellInput2[6]), .B(
        Red_SignaltoCheck[150]), .ZN(Check1_CheckInst_0_n118) );
  NAND2_X1 Check1_CheckInst_0_U118 ( .A1(Check1_CheckInst_0_n114), .A2(
        Check1_CheckInst_0_n113), .ZN(Check1_CheckInst_0_n120) );
  NOR2_X1 Check1_CheckInst_0_U117 ( .A1(Check1_CheckInst_0_n112), .A2(
        Check1_CheckInst_0_n111), .ZN(Check1_CheckInst_0_n113) );
  NAND2_X1 Check1_CheckInst_0_U116 ( .A1(Check1_CheckInst_0_n110), .A2(
        Check1_CheckInst_0_n109), .ZN(Check1_CheckInst_0_n111) );
  NOR2_X1 Check1_CheckInst_0_U115 ( .A1(Check1_CheckInst_0_n108), .A2(
        Check1_CheckInst_0_n107), .ZN(Check1_CheckInst_0_n109) );
  XOR2_X1 Check1_CheckInst_0_U114 ( .A(Red_MC_output[6]), .B(
        Red_SignaltoCheck[198]), .Z(Check1_CheckInst_0_n107) );
  XOR2_X1 Check1_CheckInst_0_U113 ( .A(Red_MC_output[12]), .B(
        Red_SignaltoCheck[204]), .Z(Check1_CheckInst_0_n108) );
  XNOR2_X1 Check1_CheckInst_0_U112 ( .A(Red_MC_output[9]), .B(
        Red_SignaltoCheck[201]), .ZN(Check1_CheckInst_0_n110) );
  NAND2_X1 Check1_CheckInst_0_U111 ( .A1(Check1_CheckInst_0_n106), .A2(
        Check1_CheckInst_0_n105), .ZN(Check1_CheckInst_0_n112) );
  NOR2_X1 Check1_CheckInst_0_U110 ( .A1(Check1_CheckInst_0_n104), .A2(
        Check1_CheckInst_0_n103), .ZN(Check1_CheckInst_0_n105) );
  NAND2_X1 Check1_CheckInst_0_U109 ( .A1(Check1_CheckInst_0_n102), .A2(
        Check1_CheckInst_0_n101), .ZN(Check1_CheckInst_0_n103) );
  NOR2_X1 Check1_CheckInst_0_U108 ( .A1(Check1_CheckInst_0_n100), .A2(
        Check1_CheckInst_0_n99), .ZN(Check1_CheckInst_0_n101) );
  XOR2_X1 Check1_CheckInst_0_U107 ( .A(Red_SubCellInput2[33]), .B(
        Red_SignaltoCheck[177]), .Z(Check1_CheckInst_0_n99) );
  XOR2_X1 Check1_CheckInst_0_U106 ( .A(Red_SubCellInput2[39]), .B(
        Red_SignaltoCheck[183]), .Z(Check1_CheckInst_0_n100) );
  XNOR2_X1 Check1_CheckInst_0_U105 ( .A(Red_MC_output[15]), .B(
        Red_SignaltoCheck[207]), .ZN(Check1_CheckInst_0_n102) );
  NAND2_X1 Check1_CheckInst_0_U104 ( .A1(Check1_CheckInst_0_n98), .A2(
        Check1_CheckInst_0_n97), .ZN(Check1_CheckInst_0_n104) );
  NOR2_X1 Check1_CheckInst_0_U103 ( .A1(Check1_CheckInst_0_n96), .A2(
        Check1_CheckInst_0_n95), .ZN(Check1_CheckInst_0_n97) );
  XOR2_X1 Check1_CheckInst_0_U102 ( .A(Red_SubCellInput2[36]), .B(
        Red_SignaltoCheck[180]), .Z(Check1_CheckInst_0_n95) );
  XOR2_X1 Check1_CheckInst_0_U101 ( .A(Red_SubCellInput2[42]), .B(
        Red_SignaltoCheck[186]), .Z(Check1_CheckInst_0_n96) );
  NOR2_X1 Check1_CheckInst_0_U100 ( .A1(Check1_CheckInst_0_n94), .A2(
        Check1_CheckInst_0_n93), .ZN(Check1_CheckInst_0_n98) );
  XOR2_X1 Check1_CheckInst_0_U99 ( .A(Red_MC_output[0]), .B(
        Red_SignaltoCheck[192]), .Z(Check1_CheckInst_0_n93) );
  XOR2_X1 Check1_CheckInst_0_U98 ( .A(Red_SubCellInput2[45]), .B(
        Red_SignaltoCheck[189]), .Z(Check1_CheckInst_0_n94) );
  XNOR2_X1 Check1_CheckInst_0_U97 ( .A(Red_SignaltoCheck[210]), .B(
        Red_MC_output[18]), .ZN(Check1_CheckInst_0_n106) );
  XNOR2_X1 Check1_CheckInst_0_U96 ( .A(Red_SignaltoCheck[195]), .B(
        Red_MC_output[3]), .ZN(Check1_CheckInst_0_n114) );
  XNOR2_X1 Check1_CheckInst_0_U95 ( .A(Red_SignaltoCheck[144]), .B(
        Red_SubCellInput2[0]), .ZN(Check1_CheckInst_0_n122) );
  NOR2_X1 Check1_CheckInst_0_U94 ( .A1(Check1_CheckInst_0_n92), .A2(
        Check1_CheckInst_0_n91), .ZN(Check1_CheckInst_0_n188) );
  NAND2_X1 Check1_CheckInst_0_U93 ( .A1(Check1_CheckInst_0_n90), .A2(
        Check1_CheckInst_0_n89), .ZN(Check1_CheckInst_0_n91) );
  NOR2_X1 Check1_CheckInst_0_U92 ( .A1(Check1_CheckInst_0_n88), .A2(
        Check1_CheckInst_0_n87), .ZN(Check1_CheckInst_0_n89) );
  NAND2_X1 Check1_CheckInst_0_U91 ( .A1(Check1_CheckInst_0_n86), .A2(
        Check1_CheckInst_0_n85), .ZN(Check1_CheckInst_0_n87) );
  NOR2_X1 Check1_CheckInst_0_U90 ( .A1(Check1_CheckInst_0_n84), .A2(
        Check1_CheckInst_0_n83), .ZN(Check1_CheckInst_0_n85) );
  NAND2_X1 Check1_CheckInst_0_U89 ( .A1(Check1_CheckInst_0_n82), .A2(
        Check1_CheckInst_0_n81), .ZN(Check1_CheckInst_0_n83) );
  NOR2_X1 Check1_CheckInst_0_U88 ( .A1(Check1_CheckInst_0_n80), .A2(
        Check1_CheckInst_0_n79), .ZN(Check1_CheckInst_0_n81) );
  XOR2_X1 Check1_CheckInst_0_U87 ( .A(Red_ShiftRowsOutput2[36]), .B(
        Red_SignaltoCheck[132]), .Z(Check1_CheckInst_0_n79) );
  XOR2_X1 Check1_CheckInst_0_U86 ( .A(Red_ShiftRowsOutput2[42]), .B(
        Red_SignaltoCheck[138]), .Z(Check1_CheckInst_0_n80) );
  NOR2_X1 Check1_CheckInst_0_U85 ( .A1(Check1_CheckInst_0_n78), .A2(
        Check1_CheckInst_0_n77), .ZN(Check1_CheckInst_0_n82) );
  XOR2_X1 Check1_CheckInst_0_U84 ( .A(Red_ShiftRowsOutput2[15]), .B(
        Red_SignaltoCheck[111]), .Z(Check1_CheckInst_0_n77) );
  XOR2_X1 Check1_CheckInst_0_U83 ( .A(Red_ShiftRowsOutput2[12]), .B(
        Red_SignaltoCheck[108]), .Z(Check1_CheckInst_0_n78) );
  NAND2_X1 Check1_CheckInst_0_U82 ( .A1(Check1_CheckInst_0_n76), .A2(
        Check1_CheckInst_0_n75), .ZN(Check1_CheckInst_0_n84) );
  XNOR2_X1 Check1_CheckInst_0_U81 ( .A(Red_ShiftRowsOutput2[21]), .B(
        Red_SignaltoCheck[117]), .ZN(Check1_CheckInst_0_n75) );
  XNOR2_X1 Check1_CheckInst_0_U80 ( .A(Red_ShiftRowsOutput2[9]), .B(
        Red_SignaltoCheck[105]), .ZN(Check1_CheckInst_0_n76) );
  NOR2_X1 Check1_CheckInst_0_U79 ( .A1(Check1_CheckInst_0_n74), .A2(
        Check1_CheckInst_0_n73), .ZN(Check1_CheckInst_0_n86) );
  XOR2_X1 Check1_CheckInst_0_U78 ( .A(Red_ShiftRowsOutput2[18]), .B(
        Red_SignaltoCheck[114]), .Z(Check1_CheckInst_0_n73) );
  XOR2_X1 Check1_CheckInst_0_U77 ( .A(Red_ShiftRowsOutput2[24]), .B(
        Red_SignaltoCheck[120]), .Z(Check1_CheckInst_0_n74) );
  NAND2_X1 Check1_CheckInst_0_U76 ( .A1(Check1_CheckInst_0_n72), .A2(
        Check1_CheckInst_0_n71), .ZN(Check1_CheckInst_0_n88) );
  NOR2_X1 Check1_CheckInst_0_U75 ( .A1(Check1_CheckInst_0_n70), .A2(
        Check1_CheckInst_0_n69), .ZN(Check1_CheckInst_0_n71) );
  NAND2_X1 Check1_CheckInst_0_U74 ( .A1(Check1_CheckInst_0_n68), .A2(
        Check1_CheckInst_0_n67), .ZN(Check1_CheckInst_0_n69) );
  NOR2_X1 Check1_CheckInst_0_U73 ( .A1(Check1_CheckInst_0_n66), .A2(
        Check1_CheckInst_0_n65), .ZN(Check1_CheckInst_0_n67) );
  XOR2_X1 Check1_CheckInst_0_U72 ( .A(Red_AddRoundKeyOutput[21]), .B(
        Red_SignaltoCheck[21]), .Z(Check1_CheckInst_0_n65) );
  XOR2_X1 Check1_CheckInst_0_U71 ( .A(Red_AddRoundKeyOutput[18]), .B(
        Red_SignaltoCheck[18]), .Z(Check1_CheckInst_0_n66) );
  NOR2_X1 Check1_CheckInst_0_U70 ( .A1(Check1_CheckInst_0_n64), .A2(
        Check1_CheckInst_0_n63), .ZN(Check1_CheckInst_0_n68) );
  XOR2_X1 Check1_CheckInst_0_U69 ( .A(Red_AddRoundKeyOutput[27]), .B(
        Red_SignaltoCheck[27]), .Z(Check1_CheckInst_0_n63) );
  XOR2_X1 Check1_CheckInst_0_U68 ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[15]), .Z(Check1_CheckInst_0_n64) );
  NAND2_X1 Check1_CheckInst_0_U67 ( .A1(Check1_CheckInst_0_n62), .A2(
        Check1_CheckInst_0_n61), .ZN(Check1_CheckInst_0_n70) );
  XNOR2_X1 Check1_CheckInst_0_U66 ( .A(Red_AddRoundKeyOutput[24]), .B(
        Red_SignaltoCheck[24]), .ZN(Check1_CheckInst_0_n61) );
  XNOR2_X1 Check1_CheckInst_0_U65 ( .A(Red_AddRoundKeyOutput[30]), .B(
        Red_SignaltoCheck[30]), .ZN(Check1_CheckInst_0_n62) );
  NOR2_X1 Check1_CheckInst_0_U64 ( .A1(Check1_CheckInst_0_n60), .A2(
        Check1_CheckInst_0_n59), .ZN(Check1_CheckInst_0_n72) );
  XOR2_X1 Check1_CheckInst_0_U63 ( .A(Red_ShiftRowsOutput[45]), .B(
        Red_SignaltoCheck[285]), .Z(Check1_CheckInst_0_n59) );
  XOR2_X1 Check1_CheckInst_0_U62 ( .A(Red_SignaltoCheck[3]), .B(
        Red_AddRoundKeyOutput[3]), .Z(Check1_CheckInst_0_n60) );
  NOR2_X1 Check1_CheckInst_0_U61 ( .A1(Check1_CheckInst_0_n58), .A2(
        Check1_CheckInst_0_n57), .ZN(Check1_CheckInst_0_n90) );
  NAND2_X1 Check1_CheckInst_0_U60 ( .A1(Check1_CheckInst_0_n56), .A2(
        Check1_CheckInst_0_n55), .ZN(Check1_CheckInst_0_n57) );
  NOR2_X1 Check1_CheckInst_0_U59 ( .A1(Check1_CheckInst_0_n54), .A2(
        Check1_CheckInst_0_n53), .ZN(Check1_CheckInst_0_n55) );
  NAND2_X1 Check1_CheckInst_0_U58 ( .A1(Check1_CheckInst_0_n52), .A2(
        Check1_CheckInst_0_n51), .ZN(Check1_CheckInst_0_n53) );
  XNOR2_X1 Check1_CheckInst_0_U57 ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[9]), .ZN(Check1_CheckInst_0_n51) );
  XNOR2_X1 Check1_CheckInst_0_U56 ( .A(Red_SignaltoCheck[0]), .B(
        Red_AddRoundKeyOutput[0]), .ZN(Check1_CheckInst_0_n52) );
  NAND2_X1 Check1_CheckInst_0_U55 ( .A1(Check1_CheckInst_0_n50), .A2(
        Check1_CheckInst_0_n49), .ZN(Check1_CheckInst_0_n54) );
  XNOR2_X1 Check1_CheckInst_0_U54 ( .A(Red_AddRoundKeyOutput[6]), .B(
        Red_SignaltoCheck[6]), .ZN(Check1_CheckInst_0_n49) );
  XNOR2_X1 Check1_CheckInst_0_U53 ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[12]), .ZN(Check1_CheckInst_0_n50) );
  NOR2_X1 Check1_CheckInst_0_U52 ( .A1(Check1_CheckInst_0_n48), .A2(
        Check1_CheckInst_0_n47), .ZN(Check1_CheckInst_0_n56) );
  XOR2_X1 Check1_CheckInst_0_U51 ( .A(Red_MC_output2[9]), .B(
        Red_SignaltoCheck[57]), .Z(Check1_CheckInst_0_n47) );
  XOR2_X1 Check1_CheckInst_0_U50 ( .A(Red_MC_output2[6]), .B(
        Red_SignaltoCheck[54]), .Z(Check1_CheckInst_0_n48) );
  NAND2_X1 Check1_CheckInst_0_U49 ( .A1(Check1_CheckInst_0_n46), .A2(
        Check1_CheckInst_0_n45), .ZN(Check1_CheckInst_0_n58) );
  XNOR2_X1 Check1_CheckInst_0_U48 ( .A(Red_MC_output2[15]), .B(
        Red_SignaltoCheck[63]), .ZN(Check1_CheckInst_0_n45) );
  XNOR2_X1 Check1_CheckInst_0_U47 ( .A(Red_MC_output2[3]), .B(
        Red_SignaltoCheck[51]), .ZN(Check1_CheckInst_0_n46) );
  NAND2_X1 Check1_CheckInst_0_U46 ( .A1(Check1_CheckInst_0_n44), .A2(
        Check1_CheckInst_0_n43), .ZN(Check1_CheckInst_0_n92) );
  NOR2_X1 Check1_CheckInst_0_U45 ( .A1(Check1_CheckInst_0_n42), .A2(
        Check1_CheckInst_0_n41), .ZN(Check1_CheckInst_0_n43) );
  NAND2_X1 Check1_CheckInst_0_U44 ( .A1(Check1_CheckInst_0_n40), .A2(
        Check1_CheckInst_0_n39), .ZN(Check1_CheckInst_0_n41) );
  NOR2_X1 Check1_CheckInst_0_U43 ( .A1(Check1_CheckInst_0_n38), .A2(
        Check1_CheckInst_0_n37), .ZN(Check1_CheckInst_0_n39) );
  XOR2_X1 Check1_CheckInst_0_U42 ( .A(Red_MC_output2[12]), .B(
        Red_SignaltoCheck[60]), .Z(Check1_CheckInst_0_n37) );
  XOR2_X1 Check1_CheckInst_0_U41 ( .A(Red_MC_output2[18]), .B(
        Red_SignaltoCheck[66]), .Z(Check1_CheckInst_0_n38) );
  NOR2_X1 Check1_CheckInst_0_U40 ( .A1(Check1_CheckInst_0_n36), .A2(
        Check1_CheckInst_0_n35), .ZN(Check1_CheckInst_0_n40) );
  XOR2_X1 Check1_CheckInst_0_U39 ( .A(Red_AddRoundKeyOutput[39]), .B(
        Red_SignaltoCheck[39]), .Z(Check1_CheckInst_0_n35) );
  XOR2_X1 Check1_CheckInst_0_U38 ( .A(Red_AddRoundKeyOutput[36]), .B(
        Red_SignaltoCheck[36]), .Z(Check1_CheckInst_0_n36) );
  NAND2_X1 Check1_CheckInst_0_U37 ( .A1(Check1_CheckInst_0_n34), .A2(
        Check1_CheckInst_0_n33), .ZN(Check1_CheckInst_0_n42) );
  XNOR2_X1 Check1_CheckInst_0_U36 ( .A(Red_AddRoundKeyOutput[45]), .B(
        Red_SignaltoCheck[45]), .ZN(Check1_CheckInst_0_n33) );
  XNOR2_X1 Check1_CheckInst_0_U35 ( .A(Red_AddRoundKeyOutput[33]), .B(
        Red_SignaltoCheck[33]), .ZN(Check1_CheckInst_0_n34) );
  NOR2_X1 Check1_CheckInst_0_U34 ( .A1(Check1_CheckInst_0_n32), .A2(
        Check1_CheckInst_0_n31), .ZN(Check1_CheckInst_0_n44) );
  XOR2_X1 Check1_CheckInst_0_U33 ( .A(Red_AddRoundKeyOutput[42]), .B(
        Red_SignaltoCheck[42]), .Z(Check1_CheckInst_0_n31) );
  XOR2_X1 Check1_CheckInst_0_U32 ( .A(Red_MC_output2[0]), .B(
        Red_SignaltoCheck[48]), .Z(Check1_CheckInst_0_n32) );
  NAND2_X1 Check1_CheckInst_0_U31 ( .A1(Check1_CheckInst_0_n30), .A2(
        Check1_CheckInst_0_n29), .ZN(Check1_CheckInst_0_n190) );
  NOR2_X1 Check1_CheckInst_0_U30 ( .A1(Check1_CheckInst_0_n28), .A2(
        Check1_CheckInst_0_n27), .ZN(Check1_CheckInst_0_n29) );
  NAND2_X1 Check1_CheckInst_0_U29 ( .A1(Check1_CheckInst_0_n26), .A2(
        Check1_CheckInst_0_n25), .ZN(Check1_CheckInst_0_n27) );
  NOR2_X1 Check1_CheckInst_0_U28 ( .A1(Check1_CheckInst_0_n24), .A2(
        Check1_CheckInst_0_n23), .ZN(Check1_CheckInst_0_n25) );
  XOR2_X1 Check1_CheckInst_0_U27 ( .A(Red_ShiftRowsOutput[9]), .B(
        Red_SignaltoCheck[249]), .Z(Check1_CheckInst_0_n23) );
  XOR2_X1 Check1_CheckInst_0_U26 ( .A(Red_ShiftRowsOutput[15]), .B(
        Red_SignaltoCheck[255]), .Z(Check1_CheckInst_0_n24) );
  XNOR2_X1 Check1_CheckInst_0_U25 ( .A(Red_ShiftRowsOutput[39]), .B(
        Red_SignaltoCheck[279]), .ZN(Check1_CheckInst_0_n26) );
  NAND2_X1 Check1_CheckInst_0_U24 ( .A1(Check1_CheckInst_0_n22), .A2(
        Check1_CheckInst_0_n21), .ZN(Check1_CheckInst_0_n28) );
  NOR2_X1 Check1_CheckInst_0_U23 ( .A1(Check1_CheckInst_0_n20), .A2(
        Check1_CheckInst_0_n19), .ZN(Check1_CheckInst_0_n21) );
  NAND2_X1 Check1_CheckInst_0_U22 ( .A1(Check1_CheckInst_0_n18), .A2(
        Check1_CheckInst_0_n17), .ZN(Check1_CheckInst_0_n19) );
  NOR2_X1 Check1_CheckInst_0_U21 ( .A1(Check1_CheckInst_0_n16), .A2(
        Check1_CheckInst_0_n15), .ZN(Check1_CheckInst_0_n17) );
  XOR2_X1 Check1_CheckInst_0_U20 ( .A(Red_ShiftRowsOutput[24]), .B(
        Red_SignaltoCheck[264]), .Z(Check1_CheckInst_0_n15) );
  XOR2_X1 Check1_CheckInst_0_U19 ( .A(Red_ShiftRowsOutput[21]), .B(
        Red_SignaltoCheck[261]), .Z(Check1_CheckInst_0_n16) );
  XNOR2_X1 Check1_CheckInst_0_U18 ( .A(Red_ShiftRowsOutput[18]), .B(
        Red_SignaltoCheck[258]), .ZN(Check1_CheckInst_0_n18) );
  NAND2_X1 Check1_CheckInst_0_U17 ( .A1(Check1_CheckInst_0_n14), .A2(
        Check1_CheckInst_0_n13), .ZN(Check1_CheckInst_0_n20) );
  NOR2_X1 Check1_CheckInst_0_U16 ( .A1(Check1_CheckInst_0_n12), .A2(
        Check1_CheckInst_0_n11), .ZN(Check1_CheckInst_0_n13) );
  NAND2_X1 Check1_CheckInst_0_U15 ( .A1(Check1_CheckInst_0_n10), .A2(
        Check1_CheckInst_0_n9), .ZN(Check1_CheckInst_0_n11) );
  NOR2_X1 Check1_CheckInst_0_U14 ( .A1(Check1_CheckInst_0_n8), .A2(
        Check1_CheckInst_0_n7), .ZN(Check1_CheckInst_0_n9) );
  XOR2_X1 Check1_CheckInst_0_U13 ( .A(Red_SubCellInput2[18]), .B(
        Red_SignaltoCheck[162]), .Z(Check1_CheckInst_0_n7) );
  XOR2_X1 Check1_CheckInst_0_U12 ( .A(Red_SubCellInput2[24]), .B(
        Red_SignaltoCheck[168]), .Z(Check1_CheckInst_0_n8) );
  XNOR2_X1 Check1_CheckInst_0_U11 ( .A(Red_SubCellInput2[21]), .B(
        Red_SignaltoCheck[165]), .ZN(Check1_CheckInst_0_n10) );
  NAND2_X1 Check1_CheckInst_0_U10 ( .A1(Check1_CheckInst_0_n6), .A2(
        Check1_CheckInst_0_n5), .ZN(Check1_CheckInst_0_n12) );
  NOR2_X1 Check1_CheckInst_0_U9 ( .A1(Check1_CheckInst_0_n4), .A2(
        Check1_CheckInst_0_n3), .ZN(Check1_CheckInst_0_n5) );
  XOR2_X1 Check1_CheckInst_0_U8 ( .A(Red_SubCellInput2[30]), .B(
        Red_SignaltoCheck[174]), .Z(Check1_CheckInst_0_n3) );
  XOR2_X1 Check1_CheckInst_0_U7 ( .A(Red_SubCellInput2[27]), .B(
        Red_SignaltoCheck[171]), .Z(Check1_CheckInst_0_n4) );
  NOR2_X1 Check1_CheckInst_0_U6 ( .A1(Check1_CheckInst_0_n2), .A2(
        Check1_CheckInst_0_n1), .ZN(Check1_CheckInst_0_n6) );
  XOR2_X1 Check1_CheckInst_0_U5 ( .A(Red_ShiftRowsOutput2[45]), .B(
        Red_SignaltoCheck[141]), .Z(Check1_CheckInst_0_n1) );
  XOR2_X1 Check1_CheckInst_0_U4 ( .A(Red_SubCellInput2[3]), .B(
        Red_SignaltoCheck[147]), .Z(Check1_CheckInst_0_n2) );
  XNOR2_X1 Check1_CheckInst_0_U3 ( .A(Red_SignaltoCheck[159]), .B(
        Red_SubCellInput2[15]), .ZN(Check1_CheckInst_0_n14) );
  XNOR2_X1 Check1_CheckInst_0_U2 ( .A(Red_SignaltoCheck[252]), .B(
        Red_ShiftRowsOutput[12]), .ZN(Check1_CheckInst_0_n22) );
  XNOR2_X1 Check1_CheckInst_0_U1 ( .A(Red_SignaltoCheck[282]), .B(
        Red_ShiftRowsOutput[42]), .ZN(Check1_CheckInst_0_n30) );
  NOR2_X1 Check1_CheckInst_1_U191 ( .A1(Check1_CheckInst_1_n192), .A2(
        Check1_CheckInst_1_n191), .ZN(Error[1]) );
  NAND2_X1 Check1_CheckInst_1_U190 ( .A1(Check1_CheckInst_1_n190), .A2(
        Check1_CheckInst_1_n189), .ZN(Check1_CheckInst_1_n191) );
  NOR2_X1 Check1_CheckInst_1_U189 ( .A1(Check1_CheckInst_1_n188), .A2(
        Check1_CheckInst_1_n187), .ZN(Check1_CheckInst_1_n189) );
  NAND2_X1 Check1_CheckInst_1_U188 ( .A1(Check1_CheckInst_1_n186), .A2(
        Check1_CheckInst_1_n185), .ZN(Check1_CheckInst_1_n187) );
  NOR2_X1 Check1_CheckInst_1_U187 ( .A1(Check1_CheckInst_1_n184), .A2(
        Check1_CheckInst_1_n183), .ZN(Check1_CheckInst_1_n185) );
  NAND2_X1 Check1_CheckInst_1_U186 ( .A1(Check1_CheckInst_1_n182), .A2(
        Check1_CheckInst_1_n181), .ZN(Check1_CheckInst_1_n183) );
  NOR2_X1 Check1_CheckInst_1_U185 ( .A1(Check1_CheckInst_1_n180), .A2(
        Check1_CheckInst_1_n179), .ZN(Check1_CheckInst_1_n181) );
  NAND2_X1 Check1_CheckInst_1_U184 ( .A1(Check1_CheckInst_1_n178), .A2(
        Check1_CheckInst_1_n177), .ZN(Check1_CheckInst_1_n179) );
  NOR2_X1 Check1_CheckInst_1_U183 ( .A1(Check1_CheckInst_1_n176), .A2(
        Check1_CheckInst_1_n175), .ZN(Check1_CheckInst_1_n177) );
  NAND2_X1 Check1_CheckInst_1_U182 ( .A1(Check1_CheckInst_1_n174), .A2(
        Check1_CheckInst_1_n173), .ZN(Check1_CheckInst_1_n175) );
  XNOR2_X1 Check1_CheckInst_1_U181 ( .A(Red_ShiftRowsOutput[31]), .B(
        Red_SignaltoCheck[271]), .ZN(Check1_CheckInst_1_n173) );
  XNOR2_X1 Check1_CheckInst_1_U180 ( .A(Red_ShiftRowsOutput[37]), .B(
        Red_SignaltoCheck[277]), .ZN(Check1_CheckInst_1_n174) );
  NAND2_X1 Check1_CheckInst_1_U179 ( .A1(Check1_CheckInst_1_n172), .A2(
        Check1_CheckInst_1_n171), .ZN(Check1_CheckInst_1_n176) );
  XNOR2_X1 Check1_CheckInst_1_U178 ( .A(Red_ShiftRowsOutput[28]), .B(
        Red_SignaltoCheck[268]), .ZN(Check1_CheckInst_1_n171) );
  XNOR2_X1 Check1_CheckInst_1_U177 ( .A(Red_ShiftRowsOutput[34]), .B(
        Red_SignaltoCheck[274]), .ZN(Check1_CheckInst_1_n172) );
  NOR2_X1 Check1_CheckInst_1_U176 ( .A1(Check1_CheckInst_1_n170), .A2(
        Check1_CheckInst_1_n169), .ZN(Check1_CheckInst_1_n178) );
  XOR2_X1 Check1_CheckInst_1_U175 ( .A(Red_MC_output[37]), .B(
        Red_SignaltoCheck[229]), .Z(Check1_CheckInst_1_n169) );
  XOR2_X1 Check1_CheckInst_1_U174 ( .A(Red_MC_output[34]), .B(
        Red_SignaltoCheck[226]), .Z(Check1_CheckInst_1_n170) );
  NAND2_X1 Check1_CheckInst_1_U173 ( .A1(Check1_CheckInst_1_n168), .A2(
        Check1_CheckInst_1_n167), .ZN(Check1_CheckInst_1_n180) );
  XNOR2_X1 Check1_CheckInst_1_U172 ( .A(Red_MC_output[25]), .B(
        Red_SignaltoCheck[217]), .ZN(Check1_CheckInst_1_n167) );
  XNOR2_X1 Check1_CheckInst_1_U171 ( .A(Red_MC_output[31]), .B(
        Red_SignaltoCheck[223]), .ZN(Check1_CheckInst_1_n168) );
  NOR2_X1 Check1_CheckInst_1_U170 ( .A1(Check1_CheckInst_1_n166), .A2(
        Check1_CheckInst_1_n165), .ZN(Check1_CheckInst_1_n182) );
  NAND2_X1 Check1_CheckInst_1_U169 ( .A1(Check1_CheckInst_1_n164), .A2(
        Check1_CheckInst_1_n163), .ZN(Check1_CheckInst_1_n165) );
  NOR2_X1 Check1_CheckInst_1_U168 ( .A1(Check1_CheckInst_1_n162), .A2(
        Check1_CheckInst_1_n161), .ZN(Check1_CheckInst_1_n163) );
  NAND2_X1 Check1_CheckInst_1_U167 ( .A1(Check1_CheckInst_1_n160), .A2(
        Check1_CheckInst_1_n159), .ZN(Check1_CheckInst_1_n161) );
  XNOR2_X1 Check1_CheckInst_1_U166 ( .A(Red_MC_output[22]), .B(
        Red_SignaltoCheck[214]), .ZN(Check1_CheckInst_1_n159) );
  XNOR2_X1 Check1_CheckInst_1_U165 ( .A(Red_MC_output[28]), .B(
        Red_SignaltoCheck[220]), .ZN(Check1_CheckInst_1_n160) );
  NAND2_X1 Check1_CheckInst_1_U164 ( .A1(Check1_CheckInst_1_n158), .A2(
        Check1_CheckInst_1_n157), .ZN(Check1_CheckInst_1_n162) );
  XNOR2_X1 Check1_CheckInst_1_U163 ( .A(Red_ShiftRowsOutput[7]), .B(
        Red_SignaltoCheck[247]), .ZN(Check1_CheckInst_1_n157) );
  XNOR2_X1 Check1_CheckInst_1_U162 ( .A(Red_ShiftRowsOutput[4]), .B(
        Red_SignaltoCheck[244]), .ZN(Check1_CheckInst_1_n158) );
  NOR2_X1 Check1_CheckInst_1_U161 ( .A1(Check1_CheckInst_1_n156), .A2(
        Check1_CheckInst_1_n155), .ZN(Check1_CheckInst_1_n164) );
  XOR2_X1 Check1_CheckInst_1_U160 ( .A(Red_MC_output[43]), .B(
        Red_SignaltoCheck[235]), .Z(Check1_CheckInst_1_n155) );
  XOR2_X1 Check1_CheckInst_1_U159 ( .A(Red_ShiftRowsOutput[1]), .B(
        Red_SignaltoCheck[241]), .Z(Check1_CheckInst_1_n156) );
  NAND2_X1 Check1_CheckInst_1_U158 ( .A1(Check1_CheckInst_1_n154), .A2(
        Check1_CheckInst_1_n153), .ZN(Check1_CheckInst_1_n166) );
  XNOR2_X1 Check1_CheckInst_1_U157 ( .A(Red_MC_output[40]), .B(
        Red_SignaltoCheck[232]), .ZN(Check1_CheckInst_1_n153) );
  XNOR2_X1 Check1_CheckInst_1_U156 ( .A(Red_MC_output[46]), .B(
        Red_SignaltoCheck[238]), .ZN(Check1_CheckInst_1_n154) );
  NAND2_X1 Check1_CheckInst_1_U155 ( .A1(Check1_CheckInst_1_n152), .A2(
        Check1_CheckInst_1_n151), .ZN(Check1_CheckInst_1_n184) );
  NOR2_X1 Check1_CheckInst_1_U154 ( .A1(Check1_CheckInst_1_n150), .A2(
        Check1_CheckInst_1_n149), .ZN(Check1_CheckInst_1_n151) );
  NAND2_X1 Check1_CheckInst_1_U153 ( .A1(Check1_CheckInst_1_n148), .A2(
        Check1_CheckInst_1_n147), .ZN(Check1_CheckInst_1_n149) );
  NOR2_X1 Check1_CheckInst_1_U152 ( .A1(Check1_CheckInst_1_n146), .A2(
        Check1_CheckInst_1_n145), .ZN(Check1_CheckInst_1_n147) );
  XOR2_X1 Check1_CheckInst_1_U151 ( .A(Red_MC_output2[46]), .B(
        Red_SignaltoCheck[94]), .Z(Check1_CheckInst_1_n145) );
  XOR2_X1 Check1_CheckInst_1_U150 ( .A(Red_MC_output2[43]), .B(
        Red_SignaltoCheck[91]), .Z(Check1_CheckInst_1_n146) );
  NOR2_X1 Check1_CheckInst_1_U149 ( .A1(Check1_CheckInst_1_n144), .A2(
        Check1_CheckInst_1_n143), .ZN(Check1_CheckInst_1_n148) );
  XOR2_X1 Check1_CheckInst_1_U148 ( .A(Red_ShiftRowsOutput2[4]), .B(
        Red_SignaltoCheck[100]), .Z(Check1_CheckInst_1_n143) );
  XOR2_X1 Check1_CheckInst_1_U147 ( .A(Red_MC_output2[40]), .B(
        Red_SignaltoCheck[88]), .Z(Check1_CheckInst_1_n144) );
  NAND2_X1 Check1_CheckInst_1_U146 ( .A1(Check1_CheckInst_1_n142), .A2(
        Check1_CheckInst_1_n141), .ZN(Check1_CheckInst_1_n150) );
  XNOR2_X1 Check1_CheckInst_1_U145 ( .A(Red_ShiftRowsOutput2[1]), .B(
        Red_SignaltoCheck[97]), .ZN(Check1_CheckInst_1_n141) );
  XNOR2_X1 Check1_CheckInst_1_U144 ( .A(Red_ShiftRowsOutput2[7]), .B(
        Red_SignaltoCheck[103]), .ZN(Check1_CheckInst_1_n142) );
  NOR2_X1 Check1_CheckInst_1_U143 ( .A1(Check1_CheckInst_1_n140), .A2(
        Check1_CheckInst_1_n139), .ZN(Check1_CheckInst_1_n152) );
  XOR2_X1 Check1_CheckInst_1_U142 ( .A(Red_MC_output2[28]), .B(
        Red_SignaltoCheck[76]), .Z(Check1_CheckInst_1_n139) );
  XOR2_X1 Check1_CheckInst_1_U141 ( .A(Red_MC_output2[25]), .B(
        Red_SignaltoCheck[73]), .Z(Check1_CheckInst_1_n140) );
  NOR2_X1 Check1_CheckInst_1_U140 ( .A1(Check1_CheckInst_1_n138), .A2(
        Check1_CheckInst_1_n137), .ZN(Check1_CheckInst_1_n186) );
  NAND2_X1 Check1_CheckInst_1_U139 ( .A1(Check1_CheckInst_1_n136), .A2(
        Check1_CheckInst_1_n135), .ZN(Check1_CheckInst_1_n137) );
  NOR2_X1 Check1_CheckInst_1_U138 ( .A1(Check1_CheckInst_1_n134), .A2(
        Check1_CheckInst_1_n133), .ZN(Check1_CheckInst_1_n135) );
  NAND2_X1 Check1_CheckInst_1_U137 ( .A1(Check1_CheckInst_1_n132), .A2(
        Check1_CheckInst_1_n131), .ZN(Check1_CheckInst_1_n133) );
  XNOR2_X1 Check1_CheckInst_1_U136 ( .A(Red_MC_output2[34]), .B(
        Red_SignaltoCheck[82]), .ZN(Check1_CheckInst_1_n131) );
  XNOR2_X1 Check1_CheckInst_1_U135 ( .A(Red_MC_output2[22]), .B(
        Red_SignaltoCheck[70]), .ZN(Check1_CheckInst_1_n132) );
  NAND2_X1 Check1_CheckInst_1_U134 ( .A1(Check1_CheckInst_1_n130), .A2(
        Check1_CheckInst_1_n129), .ZN(Check1_CheckInst_1_n134) );
  XNOR2_X1 Check1_CheckInst_1_U133 ( .A(Red_MC_output2[31]), .B(
        Red_SignaltoCheck[79]), .ZN(Check1_CheckInst_1_n129) );
  XNOR2_X1 Check1_CheckInst_1_U132 ( .A(Red_MC_output2[37]), .B(
        Red_SignaltoCheck[85]), .ZN(Check1_CheckInst_1_n130) );
  NOR2_X1 Check1_CheckInst_1_U131 ( .A1(Check1_CheckInst_1_n128), .A2(
        Check1_CheckInst_1_n127), .ZN(Check1_CheckInst_1_n136) );
  XOR2_X1 Check1_CheckInst_1_U130 ( .A(Red_ShiftRowsOutput2[34]), .B(
        Red_SignaltoCheck[130]), .Z(Check1_CheckInst_1_n127) );
  XOR2_X1 Check1_CheckInst_1_U129 ( .A(Red_ShiftRowsOutput2[31]), .B(
        Red_SignaltoCheck[127]), .Z(Check1_CheckInst_1_n128) );
  NAND2_X1 Check1_CheckInst_1_U128 ( .A1(Check1_CheckInst_1_n126), .A2(
        Check1_CheckInst_1_n125), .ZN(Check1_CheckInst_1_n138) );
  XNOR2_X1 Check1_CheckInst_1_U127 ( .A(Red_ShiftRowsOutput2[40]), .B(
        Red_SignaltoCheck[136]), .ZN(Check1_CheckInst_1_n125) );
  XNOR2_X1 Check1_CheckInst_1_U126 ( .A(Red_ShiftRowsOutput2[28]), .B(
        Red_SignaltoCheck[124]), .ZN(Check1_CheckInst_1_n126) );
  NAND2_X1 Check1_CheckInst_1_U125 ( .A1(Check1_CheckInst_1_n124), .A2(
        Check1_CheckInst_1_n123), .ZN(Check1_CheckInst_1_n188) );
  NOR2_X1 Check1_CheckInst_1_U124 ( .A1(Check1_CheckInst_1_n122), .A2(
        Check1_CheckInst_1_n121), .ZN(Check1_CheckInst_1_n123) );
  NAND2_X1 Check1_CheckInst_1_U123 ( .A1(Check1_CheckInst_1_n120), .A2(
        Check1_CheckInst_1_n119), .ZN(Check1_CheckInst_1_n121) );
  NOR2_X1 Check1_CheckInst_1_U122 ( .A1(Check1_CheckInst_1_n118), .A2(
        Check1_CheckInst_1_n117), .ZN(Check1_CheckInst_1_n119) );
  XOR2_X1 Check1_CheckInst_1_U121 ( .A(Red_SubCellInput2[13]), .B(
        Red_SignaltoCheck[157]), .Z(Check1_CheckInst_1_n117) );
  XOR2_X1 Check1_CheckInst_1_U120 ( .A(Red_SubCellInput2[10]), .B(
        Red_SignaltoCheck[154]), .Z(Check1_CheckInst_1_n118) );
  XNOR2_X1 Check1_CheckInst_1_U119 ( .A(Red_SubCellInput2[7]), .B(
        Red_SignaltoCheck[151]), .ZN(Check1_CheckInst_1_n120) );
  NAND2_X1 Check1_CheckInst_1_U118 ( .A1(Check1_CheckInst_1_n116), .A2(
        Check1_CheckInst_1_n115), .ZN(Check1_CheckInst_1_n122) );
  NOR2_X1 Check1_CheckInst_1_U117 ( .A1(Check1_CheckInst_1_n114), .A2(
        Check1_CheckInst_1_n113), .ZN(Check1_CheckInst_1_n115) );
  NAND2_X1 Check1_CheckInst_1_U116 ( .A1(Check1_CheckInst_1_n112), .A2(
        Check1_CheckInst_1_n111), .ZN(Check1_CheckInst_1_n113) );
  NOR2_X1 Check1_CheckInst_1_U115 ( .A1(Check1_CheckInst_1_n110), .A2(
        Check1_CheckInst_1_n109), .ZN(Check1_CheckInst_1_n111) );
  XOR2_X1 Check1_CheckInst_1_U114 ( .A(Red_MC_output[7]), .B(
        Red_SignaltoCheck[199]), .Z(Check1_CheckInst_1_n109) );
  XOR2_X1 Check1_CheckInst_1_U113 ( .A(Red_MC_output[13]), .B(
        Red_SignaltoCheck[205]), .Z(Check1_CheckInst_1_n110) );
  XNOR2_X1 Check1_CheckInst_1_U112 ( .A(Red_MC_output[10]), .B(
        Red_SignaltoCheck[202]), .ZN(Check1_CheckInst_1_n112) );
  NAND2_X1 Check1_CheckInst_1_U111 ( .A1(Check1_CheckInst_1_n108), .A2(
        Check1_CheckInst_1_n107), .ZN(Check1_CheckInst_1_n114) );
  NOR2_X1 Check1_CheckInst_1_U110 ( .A1(Check1_CheckInst_1_n106), .A2(
        Check1_CheckInst_1_n105), .ZN(Check1_CheckInst_1_n107) );
  NAND2_X1 Check1_CheckInst_1_U109 ( .A1(Check1_CheckInst_1_n104), .A2(
        Check1_CheckInst_1_n103), .ZN(Check1_CheckInst_1_n105) );
  NOR2_X1 Check1_CheckInst_1_U108 ( .A1(Check1_CheckInst_1_n102), .A2(
        Check1_CheckInst_1_n101), .ZN(Check1_CheckInst_1_n103) );
  XOR2_X1 Check1_CheckInst_1_U107 ( .A(Red_SubCellInput2[34]), .B(
        Red_SignaltoCheck[178]), .Z(Check1_CheckInst_1_n101) );
  XOR2_X1 Check1_CheckInst_1_U106 ( .A(Red_SubCellInput2[40]), .B(
        Red_SignaltoCheck[184]), .Z(Check1_CheckInst_1_n102) );
  XNOR2_X1 Check1_CheckInst_1_U105 ( .A(Red_MC_output[16]), .B(
        Red_SignaltoCheck[208]), .ZN(Check1_CheckInst_1_n104) );
  NAND2_X1 Check1_CheckInst_1_U104 ( .A1(Check1_CheckInst_1_n100), .A2(
        Check1_CheckInst_1_n99), .ZN(Check1_CheckInst_1_n106) );
  NOR2_X1 Check1_CheckInst_1_U103 ( .A1(Check1_CheckInst_1_n98), .A2(
        Check1_CheckInst_1_n97), .ZN(Check1_CheckInst_1_n99) );
  XOR2_X1 Check1_CheckInst_1_U102 ( .A(Red_SubCellInput2[37]), .B(
        Red_SignaltoCheck[181]), .Z(Check1_CheckInst_1_n97) );
  XOR2_X1 Check1_CheckInst_1_U101 ( .A(Red_SubCellInput2[43]), .B(
        Red_SignaltoCheck[187]), .Z(Check1_CheckInst_1_n98) );
  NOR2_X1 Check1_CheckInst_1_U100 ( .A1(Check1_CheckInst_1_n96), .A2(
        Check1_CheckInst_1_n95), .ZN(Check1_CheckInst_1_n100) );
  XOR2_X1 Check1_CheckInst_1_U99 ( .A(Red_MC_output[1]), .B(
        Red_SignaltoCheck[193]), .Z(Check1_CheckInst_1_n95) );
  XOR2_X1 Check1_CheckInst_1_U98 ( .A(Red_SubCellInput2[46]), .B(
        Red_SignaltoCheck[190]), .Z(Check1_CheckInst_1_n96) );
  XNOR2_X1 Check1_CheckInst_1_U97 ( .A(Red_SignaltoCheck[211]), .B(
        Red_MC_output[19]), .ZN(Check1_CheckInst_1_n108) );
  XNOR2_X1 Check1_CheckInst_1_U96 ( .A(Red_SignaltoCheck[196]), .B(
        Red_MC_output[4]), .ZN(Check1_CheckInst_1_n116) );
  XNOR2_X1 Check1_CheckInst_1_U95 ( .A(Red_SignaltoCheck[145]), .B(
        Red_SubCellInput2[1]), .ZN(Check1_CheckInst_1_n124) );
  NOR2_X1 Check1_CheckInst_1_U94 ( .A1(Check1_CheckInst_1_n94), .A2(
        Check1_CheckInst_1_n93), .ZN(Check1_CheckInst_1_n190) );
  NAND2_X1 Check1_CheckInst_1_U93 ( .A1(Check1_CheckInst_1_n92), .A2(
        Check1_CheckInst_1_n91), .ZN(Check1_CheckInst_1_n93) );
  NOR2_X1 Check1_CheckInst_1_U92 ( .A1(Check1_CheckInst_1_n90), .A2(
        Check1_CheckInst_1_n89), .ZN(Check1_CheckInst_1_n91) );
  NAND2_X1 Check1_CheckInst_1_U91 ( .A1(Check1_CheckInst_1_n88), .A2(
        Check1_CheckInst_1_n87), .ZN(Check1_CheckInst_1_n89) );
  NOR2_X1 Check1_CheckInst_1_U90 ( .A1(Check1_CheckInst_1_n86), .A2(
        Check1_CheckInst_1_n85), .ZN(Check1_CheckInst_1_n87) );
  NAND2_X1 Check1_CheckInst_1_U89 ( .A1(Check1_CheckInst_1_n84), .A2(
        Check1_CheckInst_1_n83), .ZN(Check1_CheckInst_1_n85) );
  NOR2_X1 Check1_CheckInst_1_U88 ( .A1(Check1_CheckInst_1_n82), .A2(
        Check1_CheckInst_1_n81), .ZN(Check1_CheckInst_1_n83) );
  XOR2_X1 Check1_CheckInst_1_U87 ( .A(Red_ShiftRowsOutput2[37]), .B(
        Red_SignaltoCheck[133]), .Z(Check1_CheckInst_1_n81) );
  XOR2_X1 Check1_CheckInst_1_U86 ( .A(Red_ShiftRowsOutput2[43]), .B(
        Red_SignaltoCheck[139]), .Z(Check1_CheckInst_1_n82) );
  NOR2_X1 Check1_CheckInst_1_U85 ( .A1(Check1_CheckInst_1_n80), .A2(
        Check1_CheckInst_1_n79), .ZN(Check1_CheckInst_1_n84) );
  XOR2_X1 Check1_CheckInst_1_U84 ( .A(Red_ShiftRowsOutput2[16]), .B(
        Red_SignaltoCheck[112]), .Z(Check1_CheckInst_1_n79) );
  XOR2_X1 Check1_CheckInst_1_U83 ( .A(Red_ShiftRowsOutput2[13]), .B(
        Red_SignaltoCheck[109]), .Z(Check1_CheckInst_1_n80) );
  NAND2_X1 Check1_CheckInst_1_U82 ( .A1(Check1_CheckInst_1_n78), .A2(
        Check1_CheckInst_1_n77), .ZN(Check1_CheckInst_1_n86) );
  XNOR2_X1 Check1_CheckInst_1_U81 ( .A(Red_ShiftRowsOutput2[22]), .B(
        Red_SignaltoCheck[118]), .ZN(Check1_CheckInst_1_n77) );
  XNOR2_X1 Check1_CheckInst_1_U80 ( .A(Red_ShiftRowsOutput2[10]), .B(
        Red_SignaltoCheck[106]), .ZN(Check1_CheckInst_1_n78) );
  NOR2_X1 Check1_CheckInst_1_U79 ( .A1(Check1_CheckInst_1_n76), .A2(
        Check1_CheckInst_1_n75), .ZN(Check1_CheckInst_1_n88) );
  XOR2_X1 Check1_CheckInst_1_U78 ( .A(Red_ShiftRowsOutput2[19]), .B(
        Red_SignaltoCheck[115]), .Z(Check1_CheckInst_1_n75) );
  XOR2_X1 Check1_CheckInst_1_U77 ( .A(Red_ShiftRowsOutput2[25]), .B(
        Red_SignaltoCheck[121]), .Z(Check1_CheckInst_1_n76) );
  NAND2_X1 Check1_CheckInst_1_U76 ( .A1(Check1_CheckInst_1_n74), .A2(
        Check1_CheckInst_1_n73), .ZN(Check1_CheckInst_1_n90) );
  NOR2_X1 Check1_CheckInst_1_U75 ( .A1(Check1_CheckInst_1_n72), .A2(
        Check1_CheckInst_1_n71), .ZN(Check1_CheckInst_1_n73) );
  NAND2_X1 Check1_CheckInst_1_U74 ( .A1(Check1_CheckInst_1_n70), .A2(
        Check1_CheckInst_1_n69), .ZN(Check1_CheckInst_1_n71) );
  NOR2_X1 Check1_CheckInst_1_U73 ( .A1(Check1_CheckInst_1_n68), .A2(
        Check1_CheckInst_1_n67), .ZN(Check1_CheckInst_1_n69) );
  XOR2_X1 Check1_CheckInst_1_U72 ( .A(Red_AddRoundKeyOutput[22]), .B(
        Red_SignaltoCheck[22]), .Z(Check1_CheckInst_1_n67) );
  XOR2_X1 Check1_CheckInst_1_U71 ( .A(Red_AddRoundKeyOutput[19]), .B(
        Red_SignaltoCheck[19]), .Z(Check1_CheckInst_1_n68) );
  NOR2_X1 Check1_CheckInst_1_U70 ( .A1(Check1_CheckInst_1_n66), .A2(
        Check1_CheckInst_1_n65), .ZN(Check1_CheckInst_1_n70) );
  XOR2_X1 Check1_CheckInst_1_U69 ( .A(Red_AddRoundKeyOutput[28]), .B(
        Red_SignaltoCheck[28]), .Z(Check1_CheckInst_1_n65) );
  XOR2_X1 Check1_CheckInst_1_U68 ( .A(Red_AddRoundKeyOutput[16]), .B(
        Red_SignaltoCheck[16]), .Z(Check1_CheckInst_1_n66) );
  NAND2_X1 Check1_CheckInst_1_U67 ( .A1(Check1_CheckInst_1_n64), .A2(
        Check1_CheckInst_1_n63), .ZN(Check1_CheckInst_1_n72) );
  XNOR2_X1 Check1_CheckInst_1_U66 ( .A(Red_AddRoundKeyOutput[25]), .B(
        Red_SignaltoCheck[25]), .ZN(Check1_CheckInst_1_n63) );
  XNOR2_X1 Check1_CheckInst_1_U65 ( .A(Red_AddRoundKeyOutput[31]), .B(
        Red_SignaltoCheck[31]), .ZN(Check1_CheckInst_1_n64) );
  NOR2_X1 Check1_CheckInst_1_U64 ( .A1(Check1_CheckInst_1_n62), .A2(
        Check1_CheckInst_1_n61), .ZN(Check1_CheckInst_1_n74) );
  XOR2_X1 Check1_CheckInst_1_U63 ( .A(Red_ShiftRowsOutput[46]), .B(
        Red_SignaltoCheck[286]), .Z(Check1_CheckInst_1_n61) );
  XOR2_X1 Check1_CheckInst_1_U62 ( .A(Red_SignaltoCheck[4]), .B(
        Red_AddRoundKeyOutput[4]), .Z(Check1_CheckInst_1_n62) );
  NOR2_X1 Check1_CheckInst_1_U61 ( .A1(Check1_CheckInst_1_n60), .A2(
        Check1_CheckInst_1_n59), .ZN(Check1_CheckInst_1_n92) );
  NAND2_X1 Check1_CheckInst_1_U60 ( .A1(Check1_CheckInst_1_n58), .A2(
        Check1_CheckInst_1_n57), .ZN(Check1_CheckInst_1_n59) );
  NOR2_X1 Check1_CheckInst_1_U59 ( .A1(Check1_CheckInst_1_n56), .A2(
        Check1_CheckInst_1_n55), .ZN(Check1_CheckInst_1_n57) );
  NAND2_X1 Check1_CheckInst_1_U58 ( .A1(Check1_CheckInst_1_n54), .A2(
        Check1_CheckInst_1_n53), .ZN(Check1_CheckInst_1_n55) );
  XNOR2_X1 Check1_CheckInst_1_U57 ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[10]), .ZN(Check1_CheckInst_1_n53) );
  XNOR2_X1 Check1_CheckInst_1_U56 ( .A(Red_SignaltoCheck[1]), .B(
        Red_AddRoundKeyOutput[1]), .ZN(Check1_CheckInst_1_n54) );
  NAND2_X1 Check1_CheckInst_1_U55 ( .A1(Check1_CheckInst_1_n52), .A2(
        Check1_CheckInst_1_n51), .ZN(Check1_CheckInst_1_n56) );
  XNOR2_X1 Check1_CheckInst_1_U54 ( .A(Red_AddRoundKeyOutput[7]), .B(
        Red_SignaltoCheck[7]), .ZN(Check1_CheckInst_1_n51) );
  XNOR2_X1 Check1_CheckInst_1_U53 ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[13]), .ZN(Check1_CheckInst_1_n52) );
  NOR2_X1 Check1_CheckInst_1_U52 ( .A1(Check1_CheckInst_1_n50), .A2(
        Check1_CheckInst_1_n49), .ZN(Check1_CheckInst_1_n58) );
  XOR2_X1 Check1_CheckInst_1_U51 ( .A(Red_MC_output2[10]), .B(
        Red_SignaltoCheck[58]), .Z(Check1_CheckInst_1_n49) );
  XOR2_X1 Check1_CheckInst_1_U50 ( .A(Red_MC_output2[7]), .B(
        Red_SignaltoCheck[55]), .Z(Check1_CheckInst_1_n50) );
  NAND2_X1 Check1_CheckInst_1_U49 ( .A1(Check1_CheckInst_1_n48), .A2(
        Check1_CheckInst_1_n47), .ZN(Check1_CheckInst_1_n60) );
  XNOR2_X1 Check1_CheckInst_1_U48 ( .A(Red_MC_output2[16]), .B(
        Red_SignaltoCheck[64]), .ZN(Check1_CheckInst_1_n47) );
  XNOR2_X1 Check1_CheckInst_1_U47 ( .A(Red_MC_output2[4]), .B(
        Red_SignaltoCheck[52]), .ZN(Check1_CheckInst_1_n48) );
  NAND2_X1 Check1_CheckInst_1_U46 ( .A1(Check1_CheckInst_1_n46), .A2(
        Check1_CheckInst_1_n45), .ZN(Check1_CheckInst_1_n94) );
  NOR2_X1 Check1_CheckInst_1_U45 ( .A1(Check1_CheckInst_1_n44), .A2(
        Check1_CheckInst_1_n43), .ZN(Check1_CheckInst_1_n45) );
  NAND2_X1 Check1_CheckInst_1_U44 ( .A1(Check1_CheckInst_1_n42), .A2(
        Check1_CheckInst_1_n41), .ZN(Check1_CheckInst_1_n43) );
  NOR2_X1 Check1_CheckInst_1_U43 ( .A1(Check1_CheckInst_1_n40), .A2(
        Check1_CheckInst_1_n39), .ZN(Check1_CheckInst_1_n41) );
  XOR2_X1 Check1_CheckInst_1_U42 ( .A(Red_MC_output2[13]), .B(
        Red_SignaltoCheck[61]), .Z(Check1_CheckInst_1_n39) );
  XOR2_X1 Check1_CheckInst_1_U41 ( .A(Red_MC_output2[19]), .B(
        Red_SignaltoCheck[67]), .Z(Check1_CheckInst_1_n40) );
  NOR2_X1 Check1_CheckInst_1_U40 ( .A1(Check1_CheckInst_1_n38), .A2(
        Check1_CheckInst_1_n37), .ZN(Check1_CheckInst_1_n42) );
  XOR2_X1 Check1_CheckInst_1_U39 ( .A(Red_AddRoundKeyOutput[40]), .B(
        Red_SignaltoCheck[40]), .Z(Check1_CheckInst_1_n37) );
  XOR2_X1 Check1_CheckInst_1_U38 ( .A(Red_AddRoundKeyOutput[37]), .B(
        Red_SignaltoCheck[37]), .Z(Check1_CheckInst_1_n38) );
  NAND2_X1 Check1_CheckInst_1_U37 ( .A1(Check1_CheckInst_1_n36), .A2(
        Check1_CheckInst_1_n35), .ZN(Check1_CheckInst_1_n44) );
  XNOR2_X1 Check1_CheckInst_1_U36 ( .A(Red_AddRoundKeyOutput[46]), .B(
        Red_SignaltoCheck[46]), .ZN(Check1_CheckInst_1_n35) );
  XNOR2_X1 Check1_CheckInst_1_U35 ( .A(Red_AddRoundKeyOutput[34]), .B(
        Red_SignaltoCheck[34]), .ZN(Check1_CheckInst_1_n36) );
  NOR2_X1 Check1_CheckInst_1_U34 ( .A1(Check1_CheckInst_1_n34), .A2(
        Check1_CheckInst_1_n33), .ZN(Check1_CheckInst_1_n46) );
  XOR2_X1 Check1_CheckInst_1_U33 ( .A(Red_AddRoundKeyOutput[43]), .B(
        Red_SignaltoCheck[43]), .Z(Check1_CheckInst_1_n33) );
  XOR2_X1 Check1_CheckInst_1_U32 ( .A(Red_MC_output2[1]), .B(
        Red_SignaltoCheck[49]), .Z(Check1_CheckInst_1_n34) );
  NAND2_X1 Check1_CheckInst_1_U31 ( .A1(Check1_CheckInst_1_n32), .A2(
        Check1_CheckInst_1_n31), .ZN(Check1_CheckInst_1_n192) );
  NOR2_X1 Check1_CheckInst_1_U30 ( .A1(Check1_CheckInst_1_n30), .A2(
        Check1_CheckInst_1_n29), .ZN(Check1_CheckInst_1_n31) );
  NAND2_X1 Check1_CheckInst_1_U29 ( .A1(Check1_CheckInst_1_n28), .A2(
        Check1_CheckInst_1_n27), .ZN(Check1_CheckInst_1_n29) );
  NOR2_X1 Check1_CheckInst_1_U28 ( .A1(Check1_CheckInst_1_n26), .A2(
        Check1_CheckInst_1_n25), .ZN(Check1_CheckInst_1_n27) );
  XOR2_X1 Check1_CheckInst_1_U27 ( .A(Red_ShiftRowsOutput[10]), .B(
        Red_SignaltoCheck[250]), .Z(Check1_CheckInst_1_n25) );
  XOR2_X1 Check1_CheckInst_1_U26 ( .A(Red_ShiftRowsOutput[16]), .B(
        Red_SignaltoCheck[256]), .Z(Check1_CheckInst_1_n26) );
  XNOR2_X1 Check1_CheckInst_1_U25 ( .A(Red_ShiftRowsOutput[40]), .B(
        Red_SignaltoCheck[280]), .ZN(Check1_CheckInst_1_n28) );
  NAND2_X1 Check1_CheckInst_1_U24 ( .A1(Check1_CheckInst_1_n24), .A2(
        Check1_CheckInst_1_n23), .ZN(Check1_CheckInst_1_n30) );
  NOR2_X1 Check1_CheckInst_1_U23 ( .A1(Check1_CheckInst_1_n22), .A2(
        Check1_CheckInst_1_n21), .ZN(Check1_CheckInst_1_n23) );
  NAND2_X1 Check1_CheckInst_1_U22 ( .A1(Check1_CheckInst_1_n20), .A2(
        Check1_CheckInst_1_n19), .ZN(Check1_CheckInst_1_n21) );
  NOR2_X1 Check1_CheckInst_1_U21 ( .A1(Check1_CheckInst_1_n18), .A2(
        Check1_CheckInst_1_n17), .ZN(Check1_CheckInst_1_n19) );
  XOR2_X1 Check1_CheckInst_1_U20 ( .A(Red_ShiftRowsOutput[25]), .B(
        Red_SignaltoCheck[265]), .Z(Check1_CheckInst_1_n17) );
  XOR2_X1 Check1_CheckInst_1_U19 ( .A(Red_ShiftRowsOutput[22]), .B(
        Red_SignaltoCheck[262]), .Z(Check1_CheckInst_1_n18) );
  XNOR2_X1 Check1_CheckInst_1_U18 ( .A(Red_ShiftRowsOutput[19]), .B(
        Red_SignaltoCheck[259]), .ZN(Check1_CheckInst_1_n20) );
  NAND2_X1 Check1_CheckInst_1_U17 ( .A1(Check1_CheckInst_1_n16), .A2(
        Check1_CheckInst_1_n15), .ZN(Check1_CheckInst_1_n22) );
  NOR2_X1 Check1_CheckInst_1_U16 ( .A1(Check1_CheckInst_1_n14), .A2(
        Check1_CheckInst_1_n13), .ZN(Check1_CheckInst_1_n15) );
  NAND2_X1 Check1_CheckInst_1_U15 ( .A1(Check1_CheckInst_1_n12), .A2(
        Check1_CheckInst_1_n11), .ZN(Check1_CheckInst_1_n13) );
  NOR2_X1 Check1_CheckInst_1_U14 ( .A1(Check1_CheckInst_1_n10), .A2(
        Check1_CheckInst_1_n9), .ZN(Check1_CheckInst_1_n11) );
  XOR2_X1 Check1_CheckInst_1_U13 ( .A(Red_SubCellInput2[19]), .B(
        Red_SignaltoCheck[163]), .Z(Check1_CheckInst_1_n9) );
  XOR2_X1 Check1_CheckInst_1_U12 ( .A(Red_SubCellInput2[25]), .B(
        Red_SignaltoCheck[169]), .Z(Check1_CheckInst_1_n10) );
  XNOR2_X1 Check1_CheckInst_1_U11 ( .A(Red_SubCellInput2[22]), .B(
        Red_SignaltoCheck[166]), .ZN(Check1_CheckInst_1_n12) );
  NAND2_X1 Check1_CheckInst_1_U10 ( .A1(Check1_CheckInst_1_n8), .A2(
        Check1_CheckInst_1_n7), .ZN(Check1_CheckInst_1_n14) );
  NOR2_X1 Check1_CheckInst_1_U9 ( .A1(Check1_CheckInst_1_n6), .A2(
        Check1_CheckInst_1_n5), .ZN(Check1_CheckInst_1_n7) );
  XOR2_X1 Check1_CheckInst_1_U8 ( .A(Red_SubCellInput2[31]), .B(
        Red_SignaltoCheck[175]), .Z(Check1_CheckInst_1_n5) );
  XOR2_X1 Check1_CheckInst_1_U7 ( .A(Red_SubCellInput2[28]), .B(
        Red_SignaltoCheck[172]), .Z(Check1_CheckInst_1_n6) );
  NOR2_X1 Check1_CheckInst_1_U6 ( .A1(Check1_CheckInst_1_n4), .A2(
        Check1_CheckInst_1_n3), .ZN(Check1_CheckInst_1_n8) );
  XOR2_X1 Check1_CheckInst_1_U5 ( .A(Red_ShiftRowsOutput2[46]), .B(
        Red_SignaltoCheck[142]), .Z(Check1_CheckInst_1_n3) );
  XOR2_X1 Check1_CheckInst_1_U4 ( .A(Red_SubCellInput2[4]), .B(
        Red_SignaltoCheck[148]), .Z(Check1_CheckInst_1_n4) );
  XNOR2_X1 Check1_CheckInst_1_U3 ( .A(Red_SignaltoCheck[160]), .B(
        Red_SubCellInput2[16]), .ZN(Check1_CheckInst_1_n16) );
  XNOR2_X1 Check1_CheckInst_1_U2 ( .A(Red_SignaltoCheck[253]), .B(
        Red_ShiftRowsOutput[13]), .ZN(Check1_CheckInst_1_n24) );
  XNOR2_X1 Check1_CheckInst_1_U1 ( .A(Red_SignaltoCheck[283]), .B(
        Red_ShiftRowsOutput[43]), .ZN(Check1_CheckInst_1_n32) );
  NOR2_X1 Check1_CheckInst_2_U191 ( .A1(Check1_CheckInst_2_n192), .A2(
        Check1_CheckInst_2_n191), .ZN(Error[2]) );
  NAND2_X1 Check1_CheckInst_2_U190 ( .A1(Check1_CheckInst_2_n190), .A2(
        Check1_CheckInst_2_n189), .ZN(Check1_CheckInst_2_n191) );
  NOR2_X1 Check1_CheckInst_2_U189 ( .A1(Check1_CheckInst_2_n188), .A2(
        Check1_CheckInst_2_n187), .ZN(Check1_CheckInst_2_n189) );
  NAND2_X1 Check1_CheckInst_2_U188 ( .A1(Check1_CheckInst_2_n186), .A2(
        Check1_CheckInst_2_n185), .ZN(Check1_CheckInst_2_n187) );
  NOR2_X1 Check1_CheckInst_2_U187 ( .A1(Check1_CheckInst_2_n184), .A2(
        Check1_CheckInst_2_n183), .ZN(Check1_CheckInst_2_n185) );
  NAND2_X1 Check1_CheckInst_2_U186 ( .A1(Check1_CheckInst_2_n182), .A2(
        Check1_CheckInst_2_n181), .ZN(Check1_CheckInst_2_n183) );
  NOR2_X1 Check1_CheckInst_2_U185 ( .A1(Check1_CheckInst_2_n180), .A2(
        Check1_CheckInst_2_n179), .ZN(Check1_CheckInst_2_n181) );
  NAND2_X1 Check1_CheckInst_2_U184 ( .A1(Check1_CheckInst_2_n178), .A2(
        Check1_CheckInst_2_n177), .ZN(Check1_CheckInst_2_n179) );
  NOR2_X1 Check1_CheckInst_2_U183 ( .A1(Check1_CheckInst_2_n176), .A2(
        Check1_CheckInst_2_n175), .ZN(Check1_CheckInst_2_n177) );
  NAND2_X1 Check1_CheckInst_2_U182 ( .A1(Check1_CheckInst_2_n174), .A2(
        Check1_CheckInst_2_n173), .ZN(Check1_CheckInst_2_n175) );
  XNOR2_X1 Check1_CheckInst_2_U181 ( .A(Red_ShiftRowsOutput[32]), .B(
        Red_SignaltoCheck[272]), .ZN(Check1_CheckInst_2_n173) );
  XNOR2_X1 Check1_CheckInst_2_U180 ( .A(Red_ShiftRowsOutput[38]), .B(
        Red_SignaltoCheck[278]), .ZN(Check1_CheckInst_2_n174) );
  NAND2_X1 Check1_CheckInst_2_U179 ( .A1(Check1_CheckInst_2_n172), .A2(
        Check1_CheckInst_2_n171), .ZN(Check1_CheckInst_2_n176) );
  XNOR2_X1 Check1_CheckInst_2_U178 ( .A(Red_ShiftRowsOutput[29]), .B(
        Red_SignaltoCheck[269]), .ZN(Check1_CheckInst_2_n171) );
  XNOR2_X1 Check1_CheckInst_2_U177 ( .A(Red_ShiftRowsOutput[35]), .B(
        Red_SignaltoCheck[275]), .ZN(Check1_CheckInst_2_n172) );
  NOR2_X1 Check1_CheckInst_2_U176 ( .A1(Check1_CheckInst_2_n170), .A2(
        Check1_CheckInst_2_n169), .ZN(Check1_CheckInst_2_n178) );
  XOR2_X1 Check1_CheckInst_2_U175 ( .A(Red_MC_output[38]), .B(
        Red_SignaltoCheck[230]), .Z(Check1_CheckInst_2_n169) );
  XOR2_X1 Check1_CheckInst_2_U174 ( .A(Red_MC_output[35]), .B(
        Red_SignaltoCheck[227]), .Z(Check1_CheckInst_2_n170) );
  NAND2_X1 Check1_CheckInst_2_U173 ( .A1(Check1_CheckInst_2_n168), .A2(
        Check1_CheckInst_2_n167), .ZN(Check1_CheckInst_2_n180) );
  XNOR2_X1 Check1_CheckInst_2_U172 ( .A(Red_MC_output[26]), .B(
        Red_SignaltoCheck[218]), .ZN(Check1_CheckInst_2_n167) );
  XNOR2_X1 Check1_CheckInst_2_U171 ( .A(Red_MC_output[32]), .B(
        Red_SignaltoCheck[224]), .ZN(Check1_CheckInst_2_n168) );
  NOR2_X1 Check1_CheckInst_2_U170 ( .A1(Check1_CheckInst_2_n166), .A2(
        Check1_CheckInst_2_n165), .ZN(Check1_CheckInst_2_n182) );
  NAND2_X1 Check1_CheckInst_2_U169 ( .A1(Check1_CheckInst_2_n164), .A2(
        Check1_CheckInst_2_n163), .ZN(Check1_CheckInst_2_n165) );
  NOR2_X1 Check1_CheckInst_2_U168 ( .A1(Check1_CheckInst_2_n162), .A2(
        Check1_CheckInst_2_n161), .ZN(Check1_CheckInst_2_n163) );
  NAND2_X1 Check1_CheckInst_2_U167 ( .A1(Check1_CheckInst_2_n160), .A2(
        Check1_CheckInst_2_n159), .ZN(Check1_CheckInst_2_n161) );
  XNOR2_X1 Check1_CheckInst_2_U166 ( .A(Red_MC_output[23]), .B(
        Red_SignaltoCheck[215]), .ZN(Check1_CheckInst_2_n159) );
  XNOR2_X1 Check1_CheckInst_2_U165 ( .A(Red_MC_output[29]), .B(
        Red_SignaltoCheck[221]), .ZN(Check1_CheckInst_2_n160) );
  NAND2_X1 Check1_CheckInst_2_U164 ( .A1(Check1_CheckInst_2_n158), .A2(
        Check1_CheckInst_2_n157), .ZN(Check1_CheckInst_2_n162) );
  XNOR2_X1 Check1_CheckInst_2_U163 ( .A(Red_ShiftRowsOutput[8]), .B(
        Red_SignaltoCheck[248]), .ZN(Check1_CheckInst_2_n157) );
  XNOR2_X1 Check1_CheckInst_2_U162 ( .A(Red_ShiftRowsOutput[5]), .B(
        Red_SignaltoCheck[245]), .ZN(Check1_CheckInst_2_n158) );
  NOR2_X1 Check1_CheckInst_2_U161 ( .A1(Check1_CheckInst_2_n156), .A2(
        Check1_CheckInst_2_n155), .ZN(Check1_CheckInst_2_n164) );
  XOR2_X1 Check1_CheckInst_2_U160 ( .A(Red_MC_output[44]), .B(
        Red_SignaltoCheck[236]), .Z(Check1_CheckInst_2_n155) );
  XOR2_X1 Check1_CheckInst_2_U159 ( .A(Red_ShiftRowsOutput[2]), .B(
        Red_SignaltoCheck[242]), .Z(Check1_CheckInst_2_n156) );
  NAND2_X1 Check1_CheckInst_2_U158 ( .A1(Check1_CheckInst_2_n154), .A2(
        Check1_CheckInst_2_n153), .ZN(Check1_CheckInst_2_n166) );
  XNOR2_X1 Check1_CheckInst_2_U157 ( .A(Red_MC_output[41]), .B(
        Red_SignaltoCheck[233]), .ZN(Check1_CheckInst_2_n153) );
  XNOR2_X1 Check1_CheckInst_2_U156 ( .A(Red_MC_output[47]), .B(
        Red_SignaltoCheck[239]), .ZN(Check1_CheckInst_2_n154) );
  NAND2_X1 Check1_CheckInst_2_U155 ( .A1(Check1_CheckInst_2_n152), .A2(
        Check1_CheckInst_2_n151), .ZN(Check1_CheckInst_2_n184) );
  NOR2_X1 Check1_CheckInst_2_U154 ( .A1(Check1_CheckInst_2_n150), .A2(
        Check1_CheckInst_2_n149), .ZN(Check1_CheckInst_2_n151) );
  NAND2_X1 Check1_CheckInst_2_U153 ( .A1(Check1_CheckInst_2_n148), .A2(
        Check1_CheckInst_2_n147), .ZN(Check1_CheckInst_2_n149) );
  NOR2_X1 Check1_CheckInst_2_U152 ( .A1(Check1_CheckInst_2_n146), .A2(
        Check1_CheckInst_2_n145), .ZN(Check1_CheckInst_2_n147) );
  XOR2_X1 Check1_CheckInst_2_U151 ( .A(Red_MC_output2[47]), .B(
        Red_SignaltoCheck[95]), .Z(Check1_CheckInst_2_n145) );
  XOR2_X1 Check1_CheckInst_2_U150 ( .A(Red_MC_output2[44]), .B(
        Red_SignaltoCheck[92]), .Z(Check1_CheckInst_2_n146) );
  NOR2_X1 Check1_CheckInst_2_U149 ( .A1(Check1_CheckInst_2_n144), .A2(
        Check1_CheckInst_2_n143), .ZN(Check1_CheckInst_2_n148) );
  XOR2_X1 Check1_CheckInst_2_U148 ( .A(Red_ShiftRowsOutput2[5]), .B(
        Red_SignaltoCheck[101]), .Z(Check1_CheckInst_2_n143) );
  XOR2_X1 Check1_CheckInst_2_U147 ( .A(Red_MC_output2[41]), .B(
        Red_SignaltoCheck[89]), .Z(Check1_CheckInst_2_n144) );
  NAND2_X1 Check1_CheckInst_2_U146 ( .A1(Check1_CheckInst_2_n142), .A2(
        Check1_CheckInst_2_n141), .ZN(Check1_CheckInst_2_n150) );
  XNOR2_X1 Check1_CheckInst_2_U145 ( .A(Red_ShiftRowsOutput2[2]), .B(
        Red_SignaltoCheck[98]), .ZN(Check1_CheckInst_2_n141) );
  XNOR2_X1 Check1_CheckInst_2_U144 ( .A(Red_ShiftRowsOutput2[8]), .B(
        Red_SignaltoCheck[104]), .ZN(Check1_CheckInst_2_n142) );
  NOR2_X1 Check1_CheckInst_2_U143 ( .A1(Check1_CheckInst_2_n140), .A2(
        Check1_CheckInst_2_n139), .ZN(Check1_CheckInst_2_n152) );
  XOR2_X1 Check1_CheckInst_2_U142 ( .A(Red_MC_output2[29]), .B(
        Red_SignaltoCheck[77]), .Z(Check1_CheckInst_2_n139) );
  XOR2_X1 Check1_CheckInst_2_U141 ( .A(Red_MC_output2[26]), .B(
        Red_SignaltoCheck[74]), .Z(Check1_CheckInst_2_n140) );
  NOR2_X1 Check1_CheckInst_2_U140 ( .A1(Check1_CheckInst_2_n138), .A2(
        Check1_CheckInst_2_n137), .ZN(Check1_CheckInst_2_n186) );
  NAND2_X1 Check1_CheckInst_2_U139 ( .A1(Check1_CheckInst_2_n136), .A2(
        Check1_CheckInst_2_n135), .ZN(Check1_CheckInst_2_n137) );
  NOR2_X1 Check1_CheckInst_2_U138 ( .A1(Check1_CheckInst_2_n134), .A2(
        Check1_CheckInst_2_n133), .ZN(Check1_CheckInst_2_n135) );
  NAND2_X1 Check1_CheckInst_2_U137 ( .A1(Check1_CheckInst_2_n132), .A2(
        Check1_CheckInst_2_n131), .ZN(Check1_CheckInst_2_n133) );
  XNOR2_X1 Check1_CheckInst_2_U136 ( .A(Red_MC_output2[35]), .B(
        Red_SignaltoCheck[83]), .ZN(Check1_CheckInst_2_n131) );
  XNOR2_X1 Check1_CheckInst_2_U135 ( .A(Red_MC_output2[23]), .B(
        Red_SignaltoCheck[71]), .ZN(Check1_CheckInst_2_n132) );
  NAND2_X1 Check1_CheckInst_2_U134 ( .A1(Check1_CheckInst_2_n130), .A2(
        Check1_CheckInst_2_n129), .ZN(Check1_CheckInst_2_n134) );
  XNOR2_X1 Check1_CheckInst_2_U133 ( .A(Red_MC_output2[32]), .B(
        Red_SignaltoCheck[80]), .ZN(Check1_CheckInst_2_n129) );
  XNOR2_X1 Check1_CheckInst_2_U132 ( .A(Red_MC_output2[38]), .B(
        Red_SignaltoCheck[86]), .ZN(Check1_CheckInst_2_n130) );
  NOR2_X1 Check1_CheckInst_2_U131 ( .A1(Check1_CheckInst_2_n128), .A2(
        Check1_CheckInst_2_n127), .ZN(Check1_CheckInst_2_n136) );
  XOR2_X1 Check1_CheckInst_2_U130 ( .A(Red_ShiftRowsOutput2[35]), .B(
        Red_SignaltoCheck[131]), .Z(Check1_CheckInst_2_n127) );
  NAND2_X1 Check1_CheckInst_2_U129 ( .A1(Check1_CheckInst_2_n126), .A2(
        Check1_CheckInst_2_n125), .ZN(Check1_CheckInst_2_n138) );
  XNOR2_X1 Check1_CheckInst_2_U128 ( .A(Red_ShiftRowsOutput2[41]), .B(
        Red_SignaltoCheck[137]), .ZN(Check1_CheckInst_2_n125) );
  XNOR2_X1 Check1_CheckInst_2_U127 ( .A(Red_ShiftRowsOutput2[29]), .B(
        Red_SignaltoCheck[125]), .ZN(Check1_CheckInst_2_n126) );
  NAND2_X1 Check1_CheckInst_2_U126 ( .A1(Check1_CheckInst_2_n124), .A2(
        Check1_CheckInst_2_n123), .ZN(Check1_CheckInst_2_n188) );
  NOR2_X1 Check1_CheckInst_2_U125 ( .A1(Check1_CheckInst_2_n122), .A2(
        Check1_CheckInst_2_n121), .ZN(Check1_CheckInst_2_n123) );
  NAND2_X1 Check1_CheckInst_2_U124 ( .A1(Check1_CheckInst_2_n120), .A2(
        Check1_CheckInst_2_n119), .ZN(Check1_CheckInst_2_n121) );
  NOR2_X1 Check1_CheckInst_2_U123 ( .A1(Check1_CheckInst_2_n118), .A2(
        Check1_CheckInst_2_n117), .ZN(Check1_CheckInst_2_n119) );
  XOR2_X1 Check1_CheckInst_2_U122 ( .A(Red_SubCellInput2[14]), .B(
        Red_SignaltoCheck[158]), .Z(Check1_CheckInst_2_n117) );
  XOR2_X1 Check1_CheckInst_2_U121 ( .A(Red_SubCellInput2[11]), .B(
        Red_SignaltoCheck[155]), .Z(Check1_CheckInst_2_n118) );
  XNOR2_X1 Check1_CheckInst_2_U120 ( .A(Red_SubCellInput2[8]), .B(
        Red_SignaltoCheck[152]), .ZN(Check1_CheckInst_2_n120) );
  NAND2_X1 Check1_CheckInst_2_U119 ( .A1(Check1_CheckInst_2_n116), .A2(
        Check1_CheckInst_2_n115), .ZN(Check1_CheckInst_2_n122) );
  NOR2_X1 Check1_CheckInst_2_U118 ( .A1(Check1_CheckInst_2_n114), .A2(
        Check1_CheckInst_2_n113), .ZN(Check1_CheckInst_2_n115) );
  NAND2_X1 Check1_CheckInst_2_U117 ( .A1(Check1_CheckInst_2_n112), .A2(
        Check1_CheckInst_2_n111), .ZN(Check1_CheckInst_2_n113) );
  NOR2_X1 Check1_CheckInst_2_U116 ( .A1(Check1_CheckInst_2_n110), .A2(
        Check1_CheckInst_2_n109), .ZN(Check1_CheckInst_2_n111) );
  XOR2_X1 Check1_CheckInst_2_U115 ( .A(Red_MC_output[8]), .B(
        Red_SignaltoCheck[200]), .Z(Check1_CheckInst_2_n109) );
  XOR2_X1 Check1_CheckInst_2_U114 ( .A(Red_MC_output[14]), .B(
        Red_SignaltoCheck[206]), .Z(Check1_CheckInst_2_n110) );
  XNOR2_X1 Check1_CheckInst_2_U113 ( .A(Red_MC_output[11]), .B(
        Red_SignaltoCheck[203]), .ZN(Check1_CheckInst_2_n112) );
  NAND2_X1 Check1_CheckInst_2_U112 ( .A1(Check1_CheckInst_2_n108), .A2(
        Check1_CheckInst_2_n107), .ZN(Check1_CheckInst_2_n114) );
  NOR2_X1 Check1_CheckInst_2_U111 ( .A1(Check1_CheckInst_2_n106), .A2(
        Check1_CheckInst_2_n105), .ZN(Check1_CheckInst_2_n107) );
  NAND2_X1 Check1_CheckInst_2_U110 ( .A1(Check1_CheckInst_2_n104), .A2(
        Check1_CheckInst_2_n103), .ZN(Check1_CheckInst_2_n105) );
  NOR2_X1 Check1_CheckInst_2_U109 ( .A1(Check1_CheckInst_2_n102), .A2(
        Check1_CheckInst_2_n101), .ZN(Check1_CheckInst_2_n103) );
  XOR2_X1 Check1_CheckInst_2_U108 ( .A(Red_SubCellInput2[35]), .B(
        Red_SignaltoCheck[179]), .Z(Check1_CheckInst_2_n101) );
  XOR2_X1 Check1_CheckInst_2_U107 ( .A(Red_SubCellInput2[41]), .B(
        Red_SignaltoCheck[185]), .Z(Check1_CheckInst_2_n102) );
  XNOR2_X1 Check1_CheckInst_2_U106 ( .A(Red_MC_output[17]), .B(
        Red_SignaltoCheck[209]), .ZN(Check1_CheckInst_2_n104) );
  NAND2_X1 Check1_CheckInst_2_U105 ( .A1(Check1_CheckInst_2_n100), .A2(
        Check1_CheckInst_2_n99), .ZN(Check1_CheckInst_2_n106) );
  NOR2_X1 Check1_CheckInst_2_U104 ( .A1(Check1_CheckInst_2_n98), .A2(
        Check1_CheckInst_2_n97), .ZN(Check1_CheckInst_2_n99) );
  XOR2_X1 Check1_CheckInst_2_U103 ( .A(Red_SubCellInput2[38]), .B(
        Red_SignaltoCheck[182]), .Z(Check1_CheckInst_2_n97) );
  XOR2_X1 Check1_CheckInst_2_U102 ( .A(Red_SubCellInput2[44]), .B(
        Red_SignaltoCheck[188]), .Z(Check1_CheckInst_2_n98) );
  NOR2_X1 Check1_CheckInst_2_U101 ( .A1(Check1_CheckInst_2_n96), .A2(
        Check1_CheckInst_2_n95), .ZN(Check1_CheckInst_2_n100) );
  XOR2_X1 Check1_CheckInst_2_U100 ( .A(Red_MC_output[2]), .B(
        Red_SignaltoCheck[194]), .Z(Check1_CheckInst_2_n95) );
  XOR2_X1 Check1_CheckInst_2_U99 ( .A(Red_SubCellInput2[47]), .B(
        Red_SignaltoCheck[191]), .Z(Check1_CheckInst_2_n96) );
  XNOR2_X1 Check1_CheckInst_2_U98 ( .A(Red_SignaltoCheck[212]), .B(
        Red_MC_output[20]), .ZN(Check1_CheckInst_2_n108) );
  XNOR2_X1 Check1_CheckInst_2_U97 ( .A(Red_SignaltoCheck[197]), .B(
        Red_MC_output[5]), .ZN(Check1_CheckInst_2_n116) );
  XNOR2_X1 Check1_CheckInst_2_U96 ( .A(Red_SignaltoCheck[146]), .B(
        Red_SubCellInput2[2]), .ZN(Check1_CheckInst_2_n124) );
  NOR2_X1 Check1_CheckInst_2_U95 ( .A1(Check1_CheckInst_2_n94), .A2(
        Check1_CheckInst_2_n93), .ZN(Check1_CheckInst_2_n190) );
  NAND2_X1 Check1_CheckInst_2_U94 ( .A1(Check1_CheckInst_2_n92), .A2(
        Check1_CheckInst_2_n91), .ZN(Check1_CheckInst_2_n93) );
  NOR2_X1 Check1_CheckInst_2_U93 ( .A1(Check1_CheckInst_2_n90), .A2(
        Check1_CheckInst_2_n89), .ZN(Check1_CheckInst_2_n91) );
  NAND2_X1 Check1_CheckInst_2_U92 ( .A1(Check1_CheckInst_2_n88), .A2(
        Check1_CheckInst_2_n87), .ZN(Check1_CheckInst_2_n89) );
  NOR2_X1 Check1_CheckInst_2_U91 ( .A1(Check1_CheckInst_2_n86), .A2(
        Check1_CheckInst_2_n85), .ZN(Check1_CheckInst_2_n87) );
  NAND2_X1 Check1_CheckInst_2_U90 ( .A1(Check1_CheckInst_2_n84), .A2(
        Check1_CheckInst_2_n83), .ZN(Check1_CheckInst_2_n85) );
  NOR2_X1 Check1_CheckInst_2_U89 ( .A1(Check1_CheckInst_2_n82), .A2(
        Check1_CheckInst_2_n81), .ZN(Check1_CheckInst_2_n83) );
  XOR2_X1 Check1_CheckInst_2_U88 ( .A(Red_ShiftRowsOutput2[38]), .B(
        Red_SignaltoCheck[134]), .Z(Check1_CheckInst_2_n81) );
  XOR2_X1 Check1_CheckInst_2_U87 ( .A(Red_ShiftRowsOutput2[44]), .B(
        Red_SignaltoCheck[140]), .Z(Check1_CheckInst_2_n82) );
  NOR2_X1 Check1_CheckInst_2_U86 ( .A1(Check1_CheckInst_2_n80), .A2(
        Check1_CheckInst_2_n79), .ZN(Check1_CheckInst_2_n84) );
  XOR2_X1 Check1_CheckInst_2_U85 ( .A(Red_ShiftRowsOutput2[17]), .B(
        Red_SignaltoCheck[113]), .Z(Check1_CheckInst_2_n79) );
  XOR2_X1 Check1_CheckInst_2_U84 ( .A(Red_ShiftRowsOutput2[14]), .B(
        Red_SignaltoCheck[110]), .Z(Check1_CheckInst_2_n80) );
  NAND2_X1 Check1_CheckInst_2_U83 ( .A1(Check1_CheckInst_2_n78), .A2(
        Check1_CheckInst_2_n77), .ZN(Check1_CheckInst_2_n86) );
  XNOR2_X1 Check1_CheckInst_2_U82 ( .A(Red_ShiftRowsOutput2[23]), .B(
        Red_SignaltoCheck[119]), .ZN(Check1_CheckInst_2_n77) );
  XNOR2_X1 Check1_CheckInst_2_U81 ( .A(Red_ShiftRowsOutput2[11]), .B(
        Red_SignaltoCheck[107]), .ZN(Check1_CheckInst_2_n78) );
  NOR2_X1 Check1_CheckInst_2_U80 ( .A1(Check1_CheckInst_2_n76), .A2(
        Check1_CheckInst_2_n75), .ZN(Check1_CheckInst_2_n88) );
  XOR2_X1 Check1_CheckInst_2_U79 ( .A(Red_ShiftRowsOutput2[26]), .B(
        Red_SignaltoCheck[122]), .Z(Check1_CheckInst_2_n76) );
  NAND2_X1 Check1_CheckInst_2_U78 ( .A1(Check1_CheckInst_2_n74), .A2(
        Check1_CheckInst_2_n73), .ZN(Check1_CheckInst_2_n90) );
  NOR2_X1 Check1_CheckInst_2_U77 ( .A1(Check1_CheckInst_2_n72), .A2(
        Check1_CheckInst_2_n71), .ZN(Check1_CheckInst_2_n73) );
  NAND2_X1 Check1_CheckInst_2_U76 ( .A1(Check1_CheckInst_2_n70), .A2(
        Check1_CheckInst_2_n69), .ZN(Check1_CheckInst_2_n71) );
  NOR2_X1 Check1_CheckInst_2_U75 ( .A1(Check1_CheckInst_2_n68), .A2(
        Check1_CheckInst_2_n67), .ZN(Check1_CheckInst_2_n69) );
  XOR2_X1 Check1_CheckInst_2_U74 ( .A(Red_AddRoundKeyOutput[23]), .B(
        Red_SignaltoCheck[23]), .Z(Check1_CheckInst_2_n67) );
  XOR2_X1 Check1_CheckInst_2_U73 ( .A(Red_AddRoundKeyOutput[20]), .B(
        Red_SignaltoCheck[20]), .Z(Check1_CheckInst_2_n68) );
  NOR2_X1 Check1_CheckInst_2_U72 ( .A1(Check1_CheckInst_2_n66), .A2(
        Check1_CheckInst_2_n65), .ZN(Check1_CheckInst_2_n70) );
  XOR2_X1 Check1_CheckInst_2_U71 ( .A(Red_AddRoundKeyOutput[29]), .B(
        Red_SignaltoCheck[29]), .Z(Check1_CheckInst_2_n65) );
  XOR2_X1 Check1_CheckInst_2_U70 ( .A(Red_AddRoundKeyOutput[17]), .B(
        Red_SignaltoCheck[17]), .Z(Check1_CheckInst_2_n66) );
  NAND2_X1 Check1_CheckInst_2_U69 ( .A1(Check1_CheckInst_2_n64), .A2(
        Check1_CheckInst_2_n63), .ZN(Check1_CheckInst_2_n72) );
  XNOR2_X1 Check1_CheckInst_2_U68 ( .A(Red_AddRoundKeyOutput[26]), .B(
        Red_SignaltoCheck[26]), .ZN(Check1_CheckInst_2_n63) );
  XNOR2_X1 Check1_CheckInst_2_U67 ( .A(Red_AddRoundKeyOutput[32]), .B(
        Red_SignaltoCheck[32]), .ZN(Check1_CheckInst_2_n64) );
  NOR2_X1 Check1_CheckInst_2_U66 ( .A1(Check1_CheckInst_2_n62), .A2(
        Check1_CheckInst_2_n61), .ZN(Check1_CheckInst_2_n74) );
  XOR2_X1 Check1_CheckInst_2_U65 ( .A(Red_SignaltoCheck[5]), .B(
        Red_AddRoundKeyOutput[5]), .Z(Check1_CheckInst_2_n62) );
  NOR2_X1 Check1_CheckInst_2_U64 ( .A1(Check1_CheckInst_2_n60), .A2(
        Check1_CheckInst_2_n59), .ZN(Check1_CheckInst_2_n92) );
  NAND2_X1 Check1_CheckInst_2_U63 ( .A1(Check1_CheckInst_2_n58), .A2(
        Check1_CheckInst_2_n57), .ZN(Check1_CheckInst_2_n59) );
  NOR2_X1 Check1_CheckInst_2_U62 ( .A1(Check1_CheckInst_2_n56), .A2(
        Check1_CheckInst_2_n55), .ZN(Check1_CheckInst_2_n57) );
  NAND2_X1 Check1_CheckInst_2_U61 ( .A1(Check1_CheckInst_2_n54), .A2(
        Check1_CheckInst_2_n53), .ZN(Check1_CheckInst_2_n55) );
  XNOR2_X1 Check1_CheckInst_2_U60 ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[11]), .ZN(Check1_CheckInst_2_n53) );
  XNOR2_X1 Check1_CheckInst_2_U59 ( .A(Red_SignaltoCheck[2]), .B(
        Red_AddRoundKeyOutput[2]), .ZN(Check1_CheckInst_2_n54) );
  NAND2_X1 Check1_CheckInst_2_U58 ( .A1(Check1_CheckInst_2_n52), .A2(
        Check1_CheckInst_2_n51), .ZN(Check1_CheckInst_2_n56) );
  XNOR2_X1 Check1_CheckInst_2_U57 ( .A(Red_AddRoundKeyOutput[8]), .B(
        Red_SignaltoCheck[8]), .ZN(Check1_CheckInst_2_n51) );
  XNOR2_X1 Check1_CheckInst_2_U56 ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[14]), .ZN(Check1_CheckInst_2_n52) );
  NOR2_X1 Check1_CheckInst_2_U55 ( .A1(Check1_CheckInst_2_n50), .A2(
        Check1_CheckInst_2_n49), .ZN(Check1_CheckInst_2_n58) );
  XOR2_X1 Check1_CheckInst_2_U54 ( .A(Red_MC_output2[11]), .B(
        Red_SignaltoCheck[59]), .Z(Check1_CheckInst_2_n49) );
  XOR2_X1 Check1_CheckInst_2_U53 ( .A(Red_MC_output2[8]), .B(
        Red_SignaltoCheck[56]), .Z(Check1_CheckInst_2_n50) );
  NAND2_X1 Check1_CheckInst_2_U52 ( .A1(Check1_CheckInst_2_n48), .A2(
        Check1_CheckInst_2_n47), .ZN(Check1_CheckInst_2_n60) );
  XNOR2_X1 Check1_CheckInst_2_U51 ( .A(Red_MC_output2[17]), .B(
        Red_SignaltoCheck[65]), .ZN(Check1_CheckInst_2_n47) );
  XNOR2_X1 Check1_CheckInst_2_U50 ( .A(Red_MC_output2[5]), .B(
        Red_SignaltoCheck[53]), .ZN(Check1_CheckInst_2_n48) );
  NAND2_X1 Check1_CheckInst_2_U49 ( .A1(Check1_CheckInst_2_n46), .A2(
        Check1_CheckInst_2_n45), .ZN(Check1_CheckInst_2_n94) );
  NOR2_X1 Check1_CheckInst_2_U48 ( .A1(Check1_CheckInst_2_n44), .A2(
        Check1_CheckInst_2_n43), .ZN(Check1_CheckInst_2_n45) );
  NAND2_X1 Check1_CheckInst_2_U47 ( .A1(Check1_CheckInst_2_n42), .A2(
        Check1_CheckInst_2_n41), .ZN(Check1_CheckInst_2_n43) );
  NOR2_X1 Check1_CheckInst_2_U46 ( .A1(Check1_CheckInst_2_n40), .A2(
        Check1_CheckInst_2_n39), .ZN(Check1_CheckInst_2_n41) );
  XOR2_X1 Check1_CheckInst_2_U45 ( .A(Red_MC_output2[14]), .B(
        Red_SignaltoCheck[62]), .Z(Check1_CheckInst_2_n39) );
  XOR2_X1 Check1_CheckInst_2_U44 ( .A(Red_MC_output2[20]), .B(
        Red_SignaltoCheck[68]), .Z(Check1_CheckInst_2_n40) );
  NOR2_X1 Check1_CheckInst_2_U43 ( .A1(Check1_CheckInst_2_n38), .A2(
        Check1_CheckInst_2_n37), .ZN(Check1_CheckInst_2_n42) );
  XOR2_X1 Check1_CheckInst_2_U42 ( .A(Red_AddRoundKeyOutput[41]), .B(
        Red_SignaltoCheck[41]), .Z(Check1_CheckInst_2_n37) );
  XOR2_X1 Check1_CheckInst_2_U41 ( .A(Red_AddRoundKeyOutput[38]), .B(
        Red_SignaltoCheck[38]), .Z(Check1_CheckInst_2_n38) );
  NAND2_X1 Check1_CheckInst_2_U40 ( .A1(Check1_CheckInst_2_n36), .A2(
        Check1_CheckInst_2_n35), .ZN(Check1_CheckInst_2_n44) );
  XNOR2_X1 Check1_CheckInst_2_U39 ( .A(Red_AddRoundKeyOutput[47]), .B(
        Red_SignaltoCheck[47]), .ZN(Check1_CheckInst_2_n35) );
  XNOR2_X1 Check1_CheckInst_2_U38 ( .A(Red_AddRoundKeyOutput[35]), .B(
        Red_SignaltoCheck[35]), .ZN(Check1_CheckInst_2_n36) );
  NOR2_X1 Check1_CheckInst_2_U37 ( .A1(Check1_CheckInst_2_n34), .A2(
        Check1_CheckInst_2_n33), .ZN(Check1_CheckInst_2_n46) );
  XOR2_X1 Check1_CheckInst_2_U36 ( .A(Red_AddRoundKeyOutput[44]), .B(
        Red_SignaltoCheck[44]), .Z(Check1_CheckInst_2_n33) );
  XOR2_X1 Check1_CheckInst_2_U35 ( .A(Red_MC_output2[2]), .B(
        Red_SignaltoCheck[50]), .Z(Check1_CheckInst_2_n34) );
  NAND2_X1 Check1_CheckInst_2_U34 ( .A1(Check1_CheckInst_2_n32), .A2(
        Check1_CheckInst_2_n31), .ZN(Check1_CheckInst_2_n192) );
  NOR2_X1 Check1_CheckInst_2_U33 ( .A1(Check1_CheckInst_2_n30), .A2(
        Check1_CheckInst_2_n29), .ZN(Check1_CheckInst_2_n31) );
  NAND2_X1 Check1_CheckInst_2_U32 ( .A1(Check1_CheckInst_2_n28), .A2(
        Check1_CheckInst_2_n27), .ZN(Check1_CheckInst_2_n29) );
  NOR2_X1 Check1_CheckInst_2_U31 ( .A1(Check1_CheckInst_2_n26), .A2(
        Check1_CheckInst_2_n25), .ZN(Check1_CheckInst_2_n27) );
  XOR2_X1 Check1_CheckInst_2_U30 ( .A(Red_ShiftRowsOutput[11]), .B(
        Red_SignaltoCheck[251]), .Z(Check1_CheckInst_2_n25) );
  XOR2_X1 Check1_CheckInst_2_U29 ( .A(Red_ShiftRowsOutput[17]), .B(
        Red_SignaltoCheck[257]), .Z(Check1_CheckInst_2_n26) );
  XNOR2_X1 Check1_CheckInst_2_U28 ( .A(Red_ShiftRowsOutput[41]), .B(
        Red_SignaltoCheck[281]), .ZN(Check1_CheckInst_2_n28) );
  NAND2_X1 Check1_CheckInst_2_U27 ( .A1(Check1_CheckInst_2_n24), .A2(
        Check1_CheckInst_2_n23), .ZN(Check1_CheckInst_2_n30) );
  NOR2_X1 Check1_CheckInst_2_U26 ( .A1(Check1_CheckInst_2_n22), .A2(
        Check1_CheckInst_2_n21), .ZN(Check1_CheckInst_2_n23) );
  NAND2_X1 Check1_CheckInst_2_U25 ( .A1(Check1_CheckInst_2_n20), .A2(
        Check1_CheckInst_2_n19), .ZN(Check1_CheckInst_2_n21) );
  NOR2_X1 Check1_CheckInst_2_U24 ( .A1(Check1_CheckInst_2_n18), .A2(
        Check1_CheckInst_2_n17), .ZN(Check1_CheckInst_2_n19) );
  XNOR2_X1 Check1_CheckInst_2_U23 ( .A(Red_ShiftRowsOutput[20]), .B(
        Red_SignaltoCheck[260]), .ZN(Check1_CheckInst_2_n20) );
  NAND2_X1 Check1_CheckInst_2_U22 ( .A1(Check1_CheckInst_2_n16), .A2(
        Check1_CheckInst_2_n15), .ZN(Check1_CheckInst_2_n22) );
  NOR2_X1 Check1_CheckInst_2_U21 ( .A1(Check1_CheckInst_2_n14), .A2(
        Check1_CheckInst_2_n13), .ZN(Check1_CheckInst_2_n15) );
  NAND2_X1 Check1_CheckInst_2_U20 ( .A1(Check1_CheckInst_2_n12), .A2(
        Check1_CheckInst_2_n11), .ZN(Check1_CheckInst_2_n13) );
  NOR2_X1 Check1_CheckInst_2_U19 ( .A1(Check1_CheckInst_2_n10), .A2(
        Check1_CheckInst_2_n9), .ZN(Check1_CheckInst_2_n11) );
  XOR2_X1 Check1_CheckInst_2_U18 ( .A(Red_SubCellInput2[20]), .B(
        Red_SignaltoCheck[164]), .Z(Check1_CheckInst_2_n9) );
  XOR2_X1 Check1_CheckInst_2_U17 ( .A(Red_SubCellInput2[26]), .B(
        Red_SignaltoCheck[170]), .Z(Check1_CheckInst_2_n10) );
  XNOR2_X1 Check1_CheckInst_2_U16 ( .A(Red_SubCellInput2[23]), .B(
        Red_SignaltoCheck[167]), .ZN(Check1_CheckInst_2_n12) );
  NAND2_X1 Check1_CheckInst_2_U15 ( .A1(Check1_CheckInst_2_n8), .A2(
        Check1_CheckInst_2_n7), .ZN(Check1_CheckInst_2_n14) );
  NOR2_X1 Check1_CheckInst_2_U14 ( .A1(Check1_CheckInst_2_n6), .A2(
        Check1_CheckInst_2_n5), .ZN(Check1_CheckInst_2_n7) );
  XOR2_X1 Check1_CheckInst_2_U13 ( .A(Red_SubCellInput2[32]), .B(
        Red_SignaltoCheck[176]), .Z(Check1_CheckInst_2_n5) );
  XOR2_X1 Check1_CheckInst_2_U12 ( .A(Red_SubCellInput2[29]), .B(
        Red_SignaltoCheck[173]), .Z(Check1_CheckInst_2_n6) );
  NOR2_X1 Check1_CheckInst_2_U11 ( .A1(Check1_CheckInst_2_n4), .A2(
        Check1_CheckInst_2_n3), .ZN(Check1_CheckInst_2_n8) );
  XOR2_X1 Check1_CheckInst_2_U10 ( .A(Red_ShiftRowsOutput2[47]), .B(
        Red_SignaltoCheck[143]), .Z(Check1_CheckInst_2_n3) );
  XOR2_X1 Check1_CheckInst_2_U9 ( .A(Red_SubCellInput2[5]), .B(
        Red_SignaltoCheck[149]), .Z(Check1_CheckInst_2_n4) );
  XNOR2_X1 Check1_CheckInst_2_U8 ( .A(Red_SignaltoCheck[161]), .B(
        Red_SubCellInput2[17]), .ZN(Check1_CheckInst_2_n16) );
  XNOR2_X1 Check1_CheckInst_2_U7 ( .A(Red_SignaltoCheck[254]), .B(
        Red_ShiftRowsOutput[14]), .ZN(Check1_CheckInst_2_n24) );
  XNOR2_X1 Check1_CheckInst_2_U6 ( .A(Red_SignaltoCheck[284]), .B(
        Red_ShiftRowsOutput[44]), .ZN(Check1_CheckInst_2_n32) );
  XOR2_X1 Check1_CheckInst_2_U5 ( .A(Red_ShiftRowsOutput[47]), .B(
        Red_SignaltoCheck[287]), .Z(Check1_CheckInst_2_n61) );
  XOR2_X1 Check1_CheckInst_2_U4 ( .A(Red_ShiftRowsOutput[23]), .B(
        Red_SignaltoCheck[263]), .Z(Check1_CheckInst_2_n18) );
  XOR2_X1 Check1_CheckInst_2_U3 ( .A(Red_ShiftRowsOutput[26]), .B(
        Red_SignaltoCheck[266]), .Z(Check1_CheckInst_2_n17) );
  XOR2_X1 Check1_CheckInst_2_U2 ( .A(Red_ShiftRowsOutput2[32]), .B(
        Red_SignaltoCheck[128]), .Z(Check1_CheckInst_2_n128) );
  XOR2_X1 Check1_CheckInst_2_U1 ( .A(Red_ShiftRowsOutput2[20]), .B(
        Red_SignaltoCheck[116]), .Z(Check1_CheckInst_2_n75) );
endmodule

